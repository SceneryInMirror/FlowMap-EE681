module kernel_2_2 ( 
    i_2_2_43_0, i_2_2_58_0, i_2_2_60_0, i_2_2_63_0, i_2_2_82_0, i_2_2_91_0,
    i_2_2_107_0, i_2_2_108_0, i_2_2_113_0, i_2_2_116_0, i_2_2_129_0,
    i_2_2_134_0, i_2_2_137_0, i_2_2_139_0, i_2_2_147_0,
    o_2_2_0_0  );
  input  i_2_2_43_0, i_2_2_58_0, i_2_2_60_0, i_2_2_63_0, i_2_2_82_0,
    i_2_2_91_0, i_2_2_107_0, i_2_2_108_0, i_2_2_113_0, i_2_2_116_0,
    i_2_2_129_0, i_2_2_134_0, i_2_2_137_0, i_2_2_139_0, i_2_2_147_0;
  output o_2_2_0_0;
  assign o_2_2_0_0 = (~i_2_2_108_0 & ((~i_2_2_113_0 & ((~i_2_2_43_0 & ((~i_2_2_60_0 & ((i_2_2_137_0 & ((~i_2_2_63_0 & ((~i_2_2_107_0 & i_2_2_129_0 & i_2_2_134_0) | (i_2_2_58_0 & i_2_2_139_0 & ~i_2_2_147_0))) | (~i_2_2_82_0 & ((i_2_2_91_0 & ((~i_2_2_116_0 & i_2_2_129_0 & ~i_2_2_139_0 & (~i_2_2_107_0 | (i_2_2_63_0 & i_2_2_147_0))) | (i_2_2_116_0 & ((i_2_2_63_0 & (~i_2_2_107_0 | ~i_2_2_147_0)) | (~i_2_2_107_0 & ~i_2_2_147_0))) | (i_2_2_58_0 & ~i_2_2_147_0))) | (~i_2_2_107_0 & ((i_2_2_58_0 & (~i_2_2_147_0 | (i_2_2_63_0 & i_2_2_129_0))) | (i_2_2_134_0 & (~i_2_2_147_0 | (i_2_2_63_0 & i_2_2_139_0))) | (i_2_2_116_0 & ((i_2_2_139_0 & ~i_2_2_147_0) | (i_2_2_63_0 & (i_2_2_129_0 | ~i_2_2_147_0)))))) | (i_2_2_58_0 & (i_2_2_116_0 | (i_2_2_63_0 & ~i_2_2_147_0))) | (i_2_2_116_0 & (i_2_2_134_0 | (i_2_2_63_0 & i_2_2_129_0 & ~i_2_2_147_0))))) | (i_2_2_58_0 & ((i_2_2_63_0 & ((i_2_2_116_0 & (~i_2_2_107_0 | ~i_2_2_147_0 | (i_2_2_91_0 & (i_2_2_129_0 | i_2_2_139_0)))) | (~i_2_2_107_0 & i_2_2_139_0))) | (i_2_2_91_0 & (i_2_2_134_0 | (~i_2_2_107_0 & i_2_2_116_0 & i_2_2_129_0))) | (~i_2_2_107_0 & (i_2_2_134_0 | (i_2_2_129_0 & ~i_2_2_147_0))) | (~i_2_2_147_0 & (i_2_2_134_0 | (i_2_2_116_0 & i_2_2_129_0))))) | (i_2_2_63_0 & ~i_2_2_107_0 & ((i_2_2_116_0 & i_2_2_134_0) | (i_2_2_129_0 & i_2_2_139_0 & ~i_2_2_147_0))) | (i_2_2_116_0 & i_2_2_134_0 & ~i_2_2_147_0))) | (i_2_2_134_0 & ((~i_2_2_147_0 & ((~i_2_2_82_0 & ((((~i_2_2_107_0 & i_2_2_139_0) | (i_2_2_91_0 & ~i_2_2_139_0)) & (i_2_2_116_0 | (i_2_2_63_0 & i_2_2_129_0))) | i_2_2_58_0 | (i_2_2_63_0 & (i_2_2_116_0 | (i_2_2_91_0 & ~i_2_2_107_0 & i_2_2_139_0))))) | (i_2_2_58_0 & (((i_2_2_63_0 | ~i_2_2_107_0) & (i_2_2_116_0 | (i_2_2_91_0 & i_2_2_129_0 & i_2_2_139_0))) | (i_2_2_139_0 & (i_2_2_116_0 | (i_2_2_63_0 & ~i_2_2_107_0))) | (i_2_2_116_0 & (~i_2_2_91_0 | i_2_2_129_0)))) | (~i_2_2_107_0 & i_2_2_116_0 & ((i_2_2_63_0 & i_2_2_139_0) | (i_2_2_91_0 & i_2_2_129_0 & ~i_2_2_139_0))))) | (i_2_2_58_0 & ((i_2_2_63_0 & (((i_2_2_129_0 | i_2_2_139_0) & ((~i_2_2_82_0 & ~i_2_2_107_0) | (i_2_2_91_0 & i_2_2_116_0))) | (~i_2_2_107_0 & i_2_2_116_0))) | (~i_2_2_82_0 & (i_2_2_116_0 | (i_2_2_91_0 & ~i_2_2_107_0 & i_2_2_129_0))) | (i_2_2_91_0 & ~i_2_2_107_0 & i_2_2_116_0 & i_2_2_139_0))) | (~i_2_2_82_0 & i_2_2_116_0 & ((i_2_2_91_0 & i_2_2_129_0 & i_2_2_139_0) | (i_2_2_63_0 & (i_2_2_129_0 | (i_2_2_91_0 & ~i_2_2_107_0))))))) | (i_2_2_58_0 & ((~i_2_2_147_0 & ((i_2_2_63_0 & ((~i_2_2_82_0 & ((i_2_2_91_0 & i_2_2_116_0) | ((i_2_2_129_0 | i_2_2_139_0) & (i_2_2_116_0 | (i_2_2_91_0 & ~i_2_2_107_0))))) | (~i_2_2_107_0 & i_2_2_116_0 & (i_2_2_91_0 | i_2_2_129_0)))) | (i_2_2_116_0 & ((~i_2_2_82_0 & (~i_2_2_107_0 | (i_2_2_91_0 & i_2_2_129_0))) | (i_2_2_129_0 & i_2_2_139_0 & i_2_2_91_0 & ~i_2_2_107_0))))) | (i_2_2_63_0 & ~i_2_2_82_0 & ~i_2_2_107_0 & i_2_2_116_0 & (i_2_2_91_0 | i_2_2_129_0 | i_2_2_139_0)))))) | (i_2_2_134_0 & ((~i_2_2_107_0 & ((i_2_2_137_0 & ((~i_2_2_147_0 & ((i_2_2_91_0 & ((i_2_2_129_0 & i_2_2_139_0) | (i_2_2_63_0 & ~i_2_2_82_0))) | (i_2_2_63_0 & i_2_2_129_0 & (i_2_2_58_0 | (~i_2_2_82_0 & i_2_2_139_0))) | (i_2_2_58_0 & (~i_2_2_82_0 | i_2_2_139_0)) | (i_2_2_116_0 & ~i_2_2_129_0))) | (i_2_2_58_0 & ~i_2_2_82_0 & (i_2_2_63_0 | (~i_2_2_129_0 & ~i_2_2_139_0) | (i_2_2_129_0 & i_2_2_139_0))))) | (~i_2_2_82_0 & ((~i_2_2_147_0 & ((i_2_2_116_0 & (i_2_2_58_0 | (i_2_2_63_0 & i_2_2_91_0 & i_2_2_139_0))) | (i_2_2_58_0 & ((i_2_2_91_0 & (i_2_2_63_0 | (i_2_2_129_0 & i_2_2_139_0))) | (i_2_2_63_0 & (i_2_2_129_0 | i_2_2_139_0)))))) | (i_2_2_58_0 & i_2_2_116_0 & (i_2_2_63_0 | (i_2_2_129_0 & (i_2_2_91_0 | i_2_2_139_0)))))) | (i_2_2_58_0 & i_2_2_116_0 & ~i_2_2_147_0 & ((i_2_2_91_0 & i_2_2_129_0) | (i_2_2_63_0 & (i_2_2_129_0 | i_2_2_139_0)))))) | (i_2_2_129_0 & ((i_2_2_91_0 & ((i_2_2_58_0 & ((~i_2_2_147_0 & ((i_2_2_63_0 & i_2_2_139_0 & (~i_2_2_82_0 | i_2_2_116_0)) | (~i_2_2_82_0 & i_2_2_116_0))) | (~i_2_2_82_0 & i_2_2_137_0 & ~i_2_2_139_0))) | (i_2_2_63_0 & ~i_2_2_116_0 & i_2_2_137_0 & ~i_2_2_139_0 & ~i_2_2_147_0))) | (i_2_2_139_0 & ((i_2_2_116_0 & ((i_2_2_58_0 & ~i_2_2_82_0 & (i_2_2_63_0 | ~i_2_2_147_0)) | (i_2_2_63_0 & i_2_2_137_0))) | (i_2_2_58_0 & ~i_2_2_82_0 & i_2_2_137_0 & ~i_2_2_147_0))))) | (i_2_2_58_0 & ((i_2_2_63_0 & ~i_2_2_82_0 & ((i_2_2_116_0 & (i_2_2_91_0 | ~i_2_2_147_0)) | (i_2_2_137_0 & (i_2_2_139_0 | ~i_2_2_147_0)))) | (i_2_2_116_0 & i_2_2_137_0 & ~i_2_2_147_0))) | (~i_2_2_82_0 & i_2_2_116_0 & i_2_2_137_0 & ~i_2_2_147_0))) | (~i_2_2_82_0 & ((~i_2_2_107_0 & ((~i_2_2_147_0 & ((i_2_2_58_0 & ((i_2_2_139_0 & ((i_2_2_63_0 & i_2_2_137_0) | (i_2_2_91_0 & i_2_2_116_0 & i_2_2_129_0))) | (i_2_2_63_0 & (i_2_2_91_0 | i_2_2_129_0) & (i_2_2_116_0 | i_2_2_137_0)) | (i_2_2_116_0 & i_2_2_137_0))) | (i_2_2_91_0 & i_2_2_116_0 & i_2_2_137_0 & i_2_2_139_0 & (i_2_2_63_0 | i_2_2_129_0)))) | (i_2_2_58_0 & i_2_2_91_0 & i_2_2_116_0 & i_2_2_129_0 & i_2_2_137_0))) | (i_2_2_58_0 & i_2_2_137_0 & ((i_2_2_63_0 & i_2_2_116_0 & (~i_2_2_91_0 | i_2_2_129_0)) | (i_2_2_91_0 & i_2_2_129_0 & ~i_2_2_134_0 & i_2_2_139_0))))) | (i_2_2_58_0 & ~i_2_2_107_0 & i_2_2_116_0 & i_2_2_137_0 & ~i_2_2_147_0 & (i_2_2_129_0 | (i_2_2_63_0 & i_2_2_91_0))))) | (~i_2_2_147_0 & ((i_2_2_116_0 & ((i_2_2_63_0 & ((~i_2_2_82_0 & ((i_2_2_60_0 & ((i_2_2_58_0 & i_2_2_91_0 & ~i_2_2_129_0 & i_2_2_137_0) | (~i_2_2_58_0 & ~i_2_2_107_0 & i_2_2_129_0 & i_2_2_134_0 & i_2_2_139_0))) | (~i_2_2_60_0 & ((i_2_2_91_0 & ((i_2_2_58_0 & i_2_2_134_0 & (~i_2_2_129_0 | i_2_2_139_0)) | (~i_2_2_58_0 & ~i_2_2_107_0 & ~i_2_2_137_0 & ((i_2_2_129_0 & ~i_2_2_139_0) | (~i_2_2_134_0 & i_2_2_139_0))))) | (i_2_2_129_0 & i_2_2_134_0 & i_2_2_58_0 & ~i_2_2_107_0))) | (i_2_2_137_0 & ((~i_2_2_91_0 & ((~i_2_2_129_0 & i_2_2_134_0) | (~i_2_2_107_0 & i_2_2_129_0 & i_2_2_139_0))) | (i_2_2_134_0 & ((~i_2_2_107_0 & i_2_2_139_0) | (i_2_2_129_0 & ~i_2_2_139_0))))) | (i_2_2_58_0 & i_2_2_91_0 & i_2_2_129_0 & ~i_2_2_134_0 & ~i_2_2_137_0 & i_2_2_139_0))) | (~i_2_2_60_0 & ((i_2_2_58_0 & ((i_2_2_91_0 & ((~i_2_2_107_0 & i_2_2_134_0 & i_2_2_137_0) | (~i_2_2_134_0 & ~i_2_2_137_0 & i_2_2_139_0 & i_2_2_107_0 & i_2_2_129_0))) | (i_2_2_129_0 & i_2_2_134_0 & i_2_2_137_0 & i_2_2_139_0))) | (~i_2_2_107_0 & i_2_2_129_0 & i_2_2_134_0 & i_2_2_137_0))) | (i_2_2_58_0 & i_2_2_60_0 & i_2_2_82_0 & i_2_2_91_0 & i_2_2_129_0 & i_2_2_137_0 & i_2_2_139_0))) | (i_2_2_58_0 & ((~i_2_2_60_0 & ((~i_2_2_82_0 & ((i_2_2_134_0 & i_2_2_137_0) | (i_2_2_91_0 & ~i_2_2_107_0 & i_2_2_129_0 & i_2_2_139_0 & (i_2_2_134_0 | i_2_2_137_0)))) | (i_2_2_91_0 & ~i_2_2_107_0 & i_2_2_129_0 & i_2_2_134_0 & i_2_2_137_0))) | (i_2_2_129_0 & i_2_2_134_0 & i_2_2_137_0 & ~i_2_2_82_0 & i_2_2_91_0 & ~i_2_2_107_0))))) | (~i_2_2_60_0 & ((~i_2_2_82_0 & ((i_2_2_63_0 & ((i_2_2_58_0 & i_2_2_129_0 & ((i_2_2_134_0 & i_2_2_137_0) | (~i_2_2_137_0 & i_2_2_139_0 & ~i_2_2_107_0 & ~i_2_2_134_0))) | (i_2_2_91_0 & ~i_2_2_116_0 & i_2_2_137_0 & (i_2_2_134_0 | (~i_2_2_107_0 & i_2_2_139_0))))) | (i_2_2_91_0 & ~i_2_2_116_0 & i_2_2_134_0 & i_2_2_137_0 & i_2_2_139_0))) | (i_2_2_91_0 & ~i_2_2_107_0 & ~i_2_2_116_0 & ~i_2_2_129_0 & i_2_2_134_0 & i_2_2_137_0 & i_2_2_139_0))))) | (~i_2_2_82_0 & i_2_2_134_0 & i_2_2_137_0 & ((~i_2_2_60_0 & ((i_2_2_139_0 & ((i_2_2_58_0 & ~i_2_2_107_0 & i_2_2_116_0) | (i_2_2_63_0 & i_2_2_91_0 & ~i_2_2_116_0 & i_2_2_129_0))) | (i_2_2_116_0 & ((i_2_2_58_0 & ~i_2_2_107_0 & (i_2_2_63_0 | (i_2_2_91_0 & i_2_2_129_0))) | (i_2_2_129_0 & ~i_2_2_139_0 & i_2_2_63_0 & i_2_2_91_0))))) | (i_2_2_58_0 & i_2_2_63_0 & i_2_2_91_0 & i_2_2_116_0 & i_2_2_129_0 & i_2_2_139_0))))) | (i_2_2_134_0 & ((~i_2_2_43_0 & ((i_2_2_137_0 & ((i_2_2_116_0 & ((i_2_2_60_0 & i_2_2_147_0 & ((i_2_2_58_0 & i_2_2_91_0 & i_2_2_107_0 & i_2_2_129_0) | (~i_2_2_107_0 & ~i_2_2_129_0 & ~i_2_2_139_0))) | (i_2_2_58_0 & ((i_2_2_63_0 & ((~i_2_2_60_0 & ~i_2_2_82_0) | (i_2_2_91_0 & ~i_2_2_107_0 & i_2_2_129_0 & ~i_2_2_139_0 & ~i_2_2_147_0))) | (~i_2_2_82_0 & ((~i_2_2_60_0 & (i_2_2_139_0 | ~i_2_2_147_0)) | (~i_2_2_91_0 & i_2_2_139_0 & ~i_2_2_147_0))))))) | (~i_2_2_107_0 & ((i_2_2_58_0 & i_2_2_139_0 & ((i_2_2_82_0 & i_2_2_91_0 & ~i_2_2_116_0 & i_2_2_129_0 & i_2_2_147_0) | (~i_2_2_60_0 & ~i_2_2_147_0))) | (~i_2_2_60_0 & ~i_2_2_82_0 & i_2_2_91_0 & ~i_2_2_116_0 & ~i_2_2_129_0 & i_2_2_147_0))) | (i_2_2_82_0 & i_2_2_91_0 & i_2_2_58_0 & i_2_2_63_0 & i_2_2_139_0 & ~i_2_2_147_0 & ~i_2_2_116_0 & i_2_2_129_0))) | (i_2_2_58_0 & i_2_2_63_0 & ((~i_2_2_107_0 & ((i_2_2_129_0 & ((~i_2_2_60_0 & ~i_2_2_147_0 & ((~i_2_2_82_0 & i_2_2_91_0 & i_2_2_116_0) | (i_2_2_82_0 & ~i_2_2_116_0 & ~i_2_2_137_0 & ~i_2_2_139_0))) | (~i_2_2_82_0 & i_2_2_91_0 & ~i_2_2_116_0 & ~i_2_2_137_0 & i_2_2_139_0 & i_2_2_147_0))) | (~i_2_2_60_0 & ~i_2_2_82_0 & i_2_2_91_0 & ~i_2_2_129_0 & ~i_2_2_139_0 & i_2_2_147_0))) | (~i_2_2_60_0 & ~i_2_2_82_0 & i_2_2_91_0 & ~i_2_2_116_0 & i_2_2_129_0 & i_2_2_139_0 & i_2_2_147_0))))) | (~i_2_2_60_0 & i_2_2_63_0 & i_2_2_137_0 & i_2_2_139_0 & ((i_2_2_107_0 & i_2_2_147_0 & i_2_2_58_0 & ~i_2_2_82_0) | (~i_2_2_58_0 & i_2_2_91_0 & ~i_2_2_107_0 & i_2_2_116_0 & i_2_2_129_0 & ~i_2_2_147_0))))) | (~i_2_2_43_0 & i_2_2_91_0 & ~i_2_2_107_0 & i_2_2_116_0 & i_2_2_137_0 & ((i_2_2_58_0 & i_2_2_63_0 & ~i_2_2_82_0 & ~i_2_2_147_0 & (i_2_2_139_0 | (~i_2_2_60_0 & i_2_2_129_0))) | (i_2_2_60_0 & i_2_2_82_0 & i_2_2_129_0 & i_2_2_139_0 & i_2_2_147_0))))) | (~i_2_2_43_0 & ((i_2_2_58_0 & ((~i_2_2_107_0 & ((i_2_2_63_0 & ((~i_2_2_82_0 & ((i_2_2_139_0 & ((i_2_2_60_0 & ((i_2_2_91_0 & i_2_2_108_0 & i_2_2_129_0 & i_2_2_137_0 & i_2_2_147_0) | (~i_2_2_91_0 & ~i_2_2_113_0 & i_2_2_116_0 & ~i_2_2_147_0))) | (i_2_2_134_0 & ~i_2_2_147_0 & ((~i_2_2_60_0 & (~i_2_2_113_0 | (i_2_2_116_0 & i_2_2_137_0))) | (~i_2_2_113_0 & i_2_2_137_0))))) | (i_2_2_91_0 & ((~i_2_2_113_0 & i_2_2_116_0 & ((~i_2_2_129_0 & i_2_2_137_0) | (~i_2_2_60_0 & ~i_2_2_147_0))) | (~i_2_2_60_0 & i_2_2_137_0 & ((~i_2_2_116_0 & ~i_2_2_129_0 & i_2_2_147_0) | (i_2_2_129_0 & i_2_2_134_0 & ~i_2_2_139_0 & ~i_2_2_147_0))))) | (~i_2_2_113_0 & i_2_2_129_0 & ~i_2_2_147_0 & ((i_2_2_134_0 & i_2_2_137_0) | (~i_2_2_60_0 & (i_2_2_116_0 | i_2_2_134_0)))))) | (~i_2_2_147_0 & ((~i_2_2_113_0 & ((i_2_2_134_0 & ((~i_2_2_60_0 & (i_2_2_116_0 | (i_2_2_91_0 & ~i_2_2_129_0 & ~i_2_2_139_0))) | (i_2_2_91_0 & i_2_2_116_0 & ~i_2_2_129_0))) | (~i_2_2_60_0 & i_2_2_91_0 & i_2_2_137_0))) | (~i_2_2_60_0 & i_2_2_82_0 & ~i_2_2_116_0 & i_2_2_137_0 & i_2_2_139_0))))) | (~i_2_2_113_0 & ((i_2_2_134_0 & ((i_2_2_137_0 & (((~i_2_2_63_0 | ~i_2_2_129_0) & (i_2_2_116_0 | (i_2_2_91_0 & ~i_2_2_147_0))) | (~i_2_2_60_0 & ~i_2_2_82_0) | (i_2_2_91_0 & i_2_2_139_0 & ~i_2_2_147_0))) | (i_2_2_116_0 & ((~i_2_2_60_0 & (~i_2_2_82_0 | (i_2_2_91_0 & i_2_2_129_0 & i_2_2_147_0))) | (i_2_2_91_0 & i_2_2_129_0 & i_2_2_139_0 & i_2_2_147_0))))) | (~i_2_2_60_0 & i_2_2_137_0 & ((i_2_2_116_0 & (i_2_2_139_0 | ~i_2_2_147_0)) | (~i_2_2_82_0 & i_2_2_91_0 & i_2_2_139_0))))) | (i_2_2_91_0 & i_2_2_108_0 & ~i_2_2_60_0 & i_2_2_82_0 & i_2_2_129_0 & i_2_2_134_0 & i_2_2_137_0 & i_2_2_139_0 & i_2_2_147_0))) | (~i_2_2_113_0 & ((i_2_2_116_0 & ((~i_2_2_60_0 & ((i_2_2_63_0 & ((i_2_2_129_0 & ((i_2_2_91_0 & i_2_2_134_0 & (i_2_2_137_0 | (i_2_2_139_0 & ~i_2_2_147_0))) | (i_2_2_137_0 & (~i_2_2_82_0 | (i_2_2_139_0 & ~i_2_2_147_0))))) | (i_2_2_134_0 & i_2_2_137_0 & i_2_2_139_0) | (~i_2_2_82_0 & ~i_2_2_147_0 & (i_2_2_134_0 | i_2_2_137_0)))) | (~i_2_2_82_0 & ((i_2_2_137_0 & i_2_2_139_0) | (i_2_2_91_0 & i_2_2_129_0 & (i_2_2_134_0 | i_2_2_139_0)))) | (i_2_2_134_0 & i_2_2_137_0 & ~i_2_2_147_0))) | (i_2_2_134_0 & ((i_2_2_129_0 & ((~i_2_2_82_0 & (i_2_2_137_0 | (i_2_2_91_0 & i_2_2_139_0 & ~i_2_2_147_0))) | (i_2_2_91_0 & i_2_2_137_0 & ~i_2_2_147_0))) | (i_2_2_137_0 & ((~i_2_2_82_0 & ~i_2_2_139_0) | (i_2_2_63_0 & i_2_2_139_0 & ~i_2_2_147_0))))) | (~i_2_2_63_0 & ~i_2_2_82_0 & i_2_2_91_0 & i_2_2_129_0 & i_2_2_137_0 & ~i_2_2_147_0))) | (~i_2_2_82_0 & i_2_2_129_0 & i_2_2_134_0 & ((~i_2_2_60_0 & (i_2_2_137_0 | (i_2_2_91_0 & i_2_2_139_0 & ~i_2_2_147_0))) | (i_2_2_137_0 & ~i_2_2_147_0 & i_2_2_63_0 & i_2_2_91_0))))) | (~i_2_2_60_0 & ~i_2_2_82_0 & ~i_2_2_116_0 & ~i_2_2_129_0 & i_2_2_139_0 & ~i_2_2_147_0 & i_2_2_134_0 & i_2_2_137_0))) | (~i_2_2_113_0 & ((i_2_2_137_0 & ((i_2_2_116_0 & ((~i_2_2_107_0 & ((i_2_2_63_0 & ((i_2_2_129_0 & ((i_2_2_91_0 & ~i_2_2_147_0 & (~i_2_2_60_0 | (~i_2_2_82_0 & ~i_2_2_139_0))) | (i_2_2_134_0 & ~i_2_2_139_0))) | (i_2_2_139_0 & ((~i_2_2_60_0 & ((i_2_2_91_0 & ~i_2_2_147_0) | (~i_2_2_82_0 & i_2_2_147_0))) | (~i_2_2_82_0 & i_2_2_134_0 & (i_2_2_91_0 | ~i_2_2_147_0)))) | (~i_2_2_60_0 & i_2_2_134_0 & ~i_2_2_147_0))) | (~i_2_2_82_0 & ~i_2_2_147_0 & ((~i_2_2_60_0 & i_2_2_129_0) | (i_2_2_91_0 & i_2_2_134_0))))) | (~i_2_2_60_0 & ((~i_2_2_82_0 & ((i_2_2_134_0 & ~i_2_2_147_0) | (i_2_2_91_0 & i_2_2_129_0 & i_2_2_139_0 & i_2_2_147_0))) | (i_2_2_91_0 & i_2_2_129_0 & i_2_2_134_0 & i_2_2_139_0 & ~i_2_2_147_0))) | (i_2_2_134_0 & i_2_2_139_0 & ~i_2_2_147_0 & ~i_2_2_82_0 & i_2_2_91_0 & i_2_2_129_0))) | (~i_2_2_60_0 & ~i_2_2_107_0 & i_2_2_134_0 & ~i_2_2_147_0 & ((i_2_2_63_0 & ~i_2_2_82_0 & i_2_2_139_0 & (i_2_2_91_0 | i_2_2_129_0)) | (i_2_2_129_0 & ~i_2_2_139_0 & (i_2_2_82_0 | i_2_2_91_0)))))) | (i_2_2_63_0 & ~i_2_2_82_0 & ~i_2_2_107_0 & i_2_2_116_0 & i_2_2_129_0 & i_2_2_134_0 & ~i_2_2_147_0 & (~i_2_2_60_0 | (~i_2_2_139_0 & (i_2_2_91_0 | i_2_2_108_0)))))))) | (~i_2_2_113_0 & ((~i_2_2_82_0 & ((~i_2_2_60_0 & ((i_2_2_58_0 & ((i_2_2_137_0 & ((~i_2_2_147_0 & ((~i_2_2_107_0 & ((i_2_2_63_0 & i_2_2_116_0 & (i_2_2_91_0 | i_2_2_129_0)) | (i_2_2_108_0 & ~i_2_2_116_0 & i_2_2_129_0 & ~i_2_2_134_0))) | (i_2_2_91_0 & i_2_2_116_0 & i_2_2_134_0 & i_2_2_139_0))) | (i_2_2_91_0 & i_2_2_107_0 & ~i_2_2_116_0 & i_2_2_134_0 & i_2_2_139_0))) | (i_2_2_91_0 & i_2_2_107_0 & i_2_2_108_0 & i_2_2_116_0 & i_2_2_134_0 & ~i_2_2_137_0 & i_2_2_139_0))) | (i_2_2_63_0 & i_2_2_91_0 & ~i_2_2_107_0 & i_2_2_108_0 & i_2_2_116_0 & ~i_2_2_129_0 & i_2_2_134_0 & ~i_2_2_137_0 & i_2_2_139_0 & ~i_2_2_147_0))) | (i_2_2_63_0 & ~i_2_2_107_0 & i_2_2_108_0 & i_2_2_116_0 & i_2_2_137_0 & ~i_2_2_139_0 & ~i_2_2_147_0 & i_2_2_129_0 & ~i_2_2_134_0))) | (i_2_2_58_0 & ~i_2_2_60_0 & i_2_2_63_0 & i_2_2_91_0 & i_2_2_129_0 & i_2_2_134_0 & i_2_2_137_0 & i_2_2_139_0 & ((~i_2_2_107_0 & i_2_2_116_0 & i_2_2_147_0) | (i_2_2_107_0 & i_2_2_108_0 & ~i_2_2_116_0 & ~i_2_2_147_0)))));
endmodule
