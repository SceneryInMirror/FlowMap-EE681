module kernel_2_5 ( 
    i_2_5_12_0, i_2_5_42_0, i_2_5_62_0, i_2_5_65_0, i_2_5_70_0, i_2_5_82_0,
    i_2_5_84_0, i_2_5_90_0, i_2_5_91_0, i_2_5_92_0, i_2_5_93_0, i_2_5_98_0,
    i_2_5_99_0, i_2_5_102_0, i_2_5_148_0,
    o_2_5_0_0  );
  input  i_2_5_12_0, i_2_5_42_0, i_2_5_62_0, i_2_5_65_0, i_2_5_70_0,
    i_2_5_82_0, i_2_5_84_0, i_2_5_90_0, i_2_5_91_0, i_2_5_92_0, i_2_5_93_0,
    i_2_5_98_0, i_2_5_99_0, i_2_5_102_0, i_2_5_148_0;
  output o_2_5_0_0;
  assign o_2_5_0_0 = (~i_2_5_92_0 & ((~i_2_5_93_0 & ((~i_2_5_98_0 & ((~i_2_5_70_0 & ((~i_2_5_90_0 & ((~i_2_5_42_0 & ((i_2_5_84_0 & ~i_2_5_99_0) | (~i_2_5_62_0 & i_2_5_65_0 & i_2_5_82_0 & i_2_5_102_0))) | (i_2_5_82_0 & ((i_2_5_12_0 & (i_2_5_148_0 | (i_2_5_62_0 & i_2_5_102_0))) | (i_2_5_42_0 & ((i_2_5_84_0 & ~i_2_5_91_0) | (i_2_5_62_0 & ~i_2_5_84_0 & ~i_2_5_148_0))) | (i_2_5_84_0 & (~i_2_5_65_0 | (i_2_5_62_0 & (i_2_5_102_0 | i_2_5_148_0)))) | (~i_2_5_91_0 & i_2_5_148_0))) | (i_2_5_42_0 & ((~i_2_5_65_0 & i_2_5_84_0) | (~i_2_5_91_0 & ~i_2_5_99_0))) | (~i_2_5_65_0 & (((~i_2_5_91_0 | (i_2_5_62_0 & i_2_5_84_0)) & (i_2_5_12_0 | i_2_5_102_0 | i_2_5_148_0)) | (i_2_5_62_0 & (~i_2_5_91_0 | ~i_2_5_99_0)) | (~i_2_5_91_0 & (i_2_5_84_0 | ~i_2_5_99_0)))) | (((i_2_5_62_0 & (~i_2_5_91_0 | ~i_2_5_99_0)) | (~i_2_5_91_0 & (i_2_5_102_0 | i_2_5_148_0))) & (i_2_5_12_0 | i_2_5_84_0)) | (~i_2_5_91_0 & (((~i_2_5_99_0 | i_2_5_148_0) & (i_2_5_62_0 | i_2_5_102_0)) | (i_2_5_12_0 & ~i_2_5_99_0))) | (i_2_5_102_0 & ((i_2_5_62_0 & ~i_2_5_99_0) | (i_2_5_84_0 & i_2_5_148_0))))) | ((i_2_5_102_0 | i_2_5_148_0) & (((i_2_5_12_0 | i_2_5_84_0) & ((~i_2_5_65_0 & (~i_2_5_91_0 | (i_2_5_62_0 & i_2_5_82_0))) | (~i_2_5_91_0 & ~i_2_5_99_0) | (i_2_5_62_0 & (i_2_5_42_0 | ~i_2_5_99_0)))) | (i_2_5_62_0 & ((~i_2_5_91_0 & ~i_2_5_99_0) | (~i_2_5_65_0 & (~i_2_5_91_0 | ~i_2_5_99_0)))) | (~i_2_5_99_0 & ((~i_2_5_65_0 & i_2_5_82_0) | (i_2_5_42_0 & ~i_2_5_91_0))))) | (i_2_5_12_0 & ((i_2_5_42_0 & ((~i_2_5_91_0 & ~i_2_5_99_0) | (i_2_5_84_0 & i_2_5_148_0) | (~i_2_5_62_0 & ~i_2_5_65_0 & i_2_5_82_0 & ~i_2_5_102_0 & ~i_2_5_148_0))) | ((~i_2_5_65_0 | ~i_2_5_91_0) & ((i_2_5_62_0 & ~i_2_5_99_0) | (i_2_5_82_0 & i_2_5_84_0))) | (~i_2_5_65_0 & ((i_2_5_84_0 & (i_2_5_102_0 | (i_2_5_62_0 & i_2_5_148_0))) | (i_2_5_62_0 & (~i_2_5_91_0 | (i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_99_0 & (~i_2_5_91_0 | i_2_5_102_0)) | (i_2_5_82_0 & i_2_5_102_0 & i_2_5_148_0))) | (i_2_5_102_0 & ((i_2_5_62_0 & ((i_2_5_84_0 & ~i_2_5_91_0) | (i_2_5_82_0 & (~i_2_5_91_0 | i_2_5_148_0)))) | (i_2_5_148_0 & (i_2_5_84_0 | ~i_2_5_91_0)))) | (i_2_5_82_0 & i_2_5_84_0 & (~i_2_5_99_0 | i_2_5_148_0)) | (i_2_5_62_0 & ~i_2_5_91_0 & i_2_5_148_0))) | ((i_2_5_62_0 | i_2_5_102_0) & ((~i_2_5_91_0 & ((i_2_5_82_0 & (~i_2_5_99_0 | (i_2_5_42_0 & i_2_5_84_0))) | (i_2_5_84_0 & i_2_5_148_0) | (~i_2_5_65_0 & ~i_2_5_99_0))) | (i_2_5_82_0 & ~i_2_5_99_0 & i_2_5_148_0))) | ((~i_2_5_91_0 | i_2_5_148_0) & ((i_2_5_42_0 & ~i_2_5_65_0 & (~i_2_5_99_0 | (i_2_5_82_0 & i_2_5_102_0))) | (i_2_5_62_0 & i_2_5_82_0 & i_2_5_84_0 & i_2_5_102_0))) | (i_2_5_62_0 & (((~i_2_5_91_0 | ~i_2_5_99_0) & ((~i_2_5_65_0 & i_2_5_84_0) | (i_2_5_42_0 & i_2_5_82_0 & i_2_5_102_0))) | (((~i_2_5_91_0 & ~i_2_5_99_0) | (~i_2_5_65_0 & i_2_5_102_0 & i_2_5_148_0)) & (i_2_5_42_0 | i_2_5_84_0)) | (~i_2_5_65_0 & i_2_5_82_0 & (~i_2_5_99_0 | (i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_91_0 & i_2_5_102_0 & i_2_5_148_0))) | (i_2_5_148_0 & ((i_2_5_102_0 & ((~i_2_5_91_0 & ~i_2_5_99_0) | (~i_2_5_65_0 & (~i_2_5_91_0 | ~i_2_5_99_0)) | (i_2_5_42_0 & ((~i_2_5_82_0 & i_2_5_84_0) | (i_2_5_82_0 & ~i_2_5_91_0))))) | (i_2_5_82_0 & ~i_2_5_91_0 & (~i_2_5_65_0 | i_2_5_84_0)))) | (~i_2_5_65_0 & i_2_5_84_0 & ~i_2_5_91_0 & ~i_2_5_99_0))) | (i_2_5_42_0 & ((i_2_5_12_0 & ((~i_2_5_82_0 & ((~i_2_5_65_0 & i_2_5_102_0 & i_2_5_148_0) | (i_2_5_62_0 & i_2_5_84_0 & ~i_2_5_90_0 & ~i_2_5_102_0 & ~i_2_5_148_0))) | (i_2_5_102_0 & ((~i_2_5_65_0 & ((~i_2_5_90_0 & ~i_2_5_91_0) | (i_2_5_82_0 & ~i_2_5_99_0))) | (i_2_5_82_0 & ((~i_2_5_91_0 & i_2_5_148_0) | (i_2_5_62_0 & ~i_2_5_99_0))) | (i_2_5_62_0 & i_2_5_84_0 & (~i_2_5_99_0 | i_2_5_148_0)))) | (i_2_5_84_0 & ((~i_2_5_65_0 & (i_2_5_82_0 | ~i_2_5_91_0)) | (~i_2_5_91_0 & i_2_5_148_0 & (i_2_5_62_0 | ~i_2_5_90_0)))) | (~i_2_5_91_0 & ((~i_2_5_99_0 & i_2_5_148_0) | (~i_2_5_90_0 & (i_2_5_82_0 | ~i_2_5_99_0)))))) | (i_2_5_82_0 & ((((~i_2_5_91_0 & i_2_5_148_0) | (~i_2_5_99_0 & i_2_5_102_0)) & ((i_2_5_84_0 & (i_2_5_62_0 | ~i_2_5_90_0)) | (i_2_5_62_0 & (~i_2_5_65_0 | ~i_2_5_90_0)))) | (i_2_5_84_0 & ((~i_2_5_65_0 & (~i_2_5_91_0 | (~i_2_5_99_0 & i_2_5_102_0))) | ((~i_2_5_90_0 | i_2_5_148_0) & ((i_2_5_62_0 & ~i_2_5_99_0) | (~i_2_5_91_0 & i_2_5_102_0))) | (i_2_5_62_0 & ~i_2_5_90_0 & ~i_2_5_91_0))) | (~i_2_5_99_0 & ((~i_2_5_65_0 & ~i_2_5_90_0) | (i_2_5_62_0 & i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_91_0 & i_2_5_102_0 & ((i_2_5_62_0 & (~i_2_5_90_0 | i_2_5_148_0)) | (~i_2_5_90_0 & i_2_5_148_0))))) | (~i_2_5_91_0 & (((~i_2_5_90_0 | i_2_5_102_0) & ((i_2_5_62_0 & (~i_2_5_99_0 | (i_2_5_84_0 & i_2_5_148_0))) | (~i_2_5_99_0 & (~i_2_5_65_0 | i_2_5_148_0)))) | ((i_2_5_62_0 | ~i_2_5_65_0) & ((~i_2_5_99_0 & i_2_5_148_0) | (i_2_5_84_0 & ~i_2_5_90_0 & i_2_5_102_0))) | (~i_2_5_65_0 & ((i_2_5_84_0 & ~i_2_5_99_0) | (i_2_5_62_0 & (~i_2_5_99_0 | (i_2_5_84_0 & i_2_5_102_0))))) | (~i_2_5_90_0 & ~i_2_5_99_0 & (i_2_5_84_0 | i_2_5_102_0)))) | (~i_2_5_65_0 & i_2_5_102_0 & i_2_5_148_0 & ((i_2_5_62_0 & (i_2_5_84_0 | ~i_2_5_90_0)) | (i_2_5_84_0 & ~i_2_5_90_0))))) | (i_2_5_148_0 & (((i_2_5_84_0 | ~i_2_5_90_0) & ((i_2_5_62_0 & ((~i_2_5_99_0 & i_2_5_102_0) | (~i_2_5_91_0 & (~i_2_5_65_0 | ~i_2_5_99_0)))) | (i_2_5_102_0 & ((~i_2_5_65_0 & (~i_2_5_91_0 | (~i_2_5_42_0 & i_2_5_82_0))) | (i_2_5_12_0 & ~i_2_5_91_0))))) | ((i_2_5_82_0 | i_2_5_102_0) & ((i_2_5_12_0 & ~i_2_5_65_0 & i_2_5_84_0) | (i_2_5_62_0 & ~i_2_5_91_0 & ~i_2_5_99_0))) | ((~i_2_5_99_0 | (i_2_5_62_0 & ~i_2_5_91_0)) & ((i_2_5_12_0 & (~i_2_5_65_0 | (i_2_5_82_0 & i_2_5_84_0))) | (i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_90_0))) | (~i_2_5_90_0 & ((i_2_5_62_0 & ((~i_2_5_65_0 & (i_2_5_12_0 | (i_2_5_84_0 & i_2_5_102_0))) | (i_2_5_12_0 & (~i_2_5_91_0 | (i_2_5_82_0 & i_2_5_102_0))) | (~i_2_5_91_0 & i_2_5_102_0) | (i_2_5_84_0 & (~i_2_5_99_0 | (i_2_5_82_0 & i_2_5_102_0))))) | (i_2_5_12_0 & ((~i_2_5_99_0 & i_2_5_102_0) | (~i_2_5_65_0 & i_2_5_70_0))) | (i_2_5_84_0 & ((~i_2_5_65_0 & (i_2_5_82_0 | ~i_2_5_91_0)) | (~i_2_5_91_0 & (~i_2_5_99_0 | i_2_5_102_0)))) | (~i_2_5_91_0 & ~i_2_5_99_0 & i_2_5_102_0))) | (i_2_5_102_0 & ((i_2_5_62_0 & ((i_2_5_12_0 & (~i_2_5_99_0 | (i_2_5_82_0 & ~i_2_5_91_0))) | (~i_2_5_65_0 & ~i_2_5_99_0) | (i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_91_0))) | (i_2_5_82_0 & ((~i_2_5_91_0 & ~i_2_5_99_0) | (~i_2_5_65_0 & (~i_2_5_91_0 | ~i_2_5_99_0)))))) | (~i_2_5_65_0 & ~i_2_5_99_0 & ((i_2_5_62_0 & (i_2_5_84_0 | ~i_2_5_91_0)) | (~i_2_5_42_0 & ~i_2_5_82_0 & i_2_5_84_0))))) | (~i_2_5_91_0 & (((i_2_5_62_0 | i_2_5_102_0) & ((~i_2_5_90_0 & ((i_2_5_12_0 & (~i_2_5_99_0 | (~i_2_5_65_0 & i_2_5_84_0))) | (~i_2_5_99_0 & (~i_2_5_65_0 | i_2_5_82_0 | i_2_5_84_0)))) | (i_2_5_12_0 & i_2_5_82_0 & ~i_2_5_99_0))) | (i_2_5_82_0 & ((~i_2_5_65_0 & ((i_2_5_62_0 & i_2_5_84_0 & ~i_2_5_90_0) | (~i_2_5_42_0 & ~i_2_5_99_0))) | (i_2_5_62_0 & ((i_2_5_84_0 & ~i_2_5_99_0) | (i_2_5_102_0 & ((i_2_5_12_0 & (i_2_5_84_0 | ~i_2_5_90_0)) | ~i_2_5_99_0 | (i_2_5_84_0 & ~i_2_5_90_0))))) | (i_2_5_12_0 & i_2_5_84_0 & ~i_2_5_90_0))) | (i_2_5_62_0 & ((i_2_5_84_0 & ((i_2_5_12_0 & (~i_2_5_99_0 | (~i_2_5_90_0 & i_2_5_102_0))) | (~i_2_5_99_0 & (~i_2_5_65_0 | i_2_5_102_0)))) | (i_2_5_102_0 & ((~i_2_5_65_0 & (~i_2_5_90_0 | ~i_2_5_99_0)) | (~i_2_5_99_0 & (i_2_5_12_0 | ~i_2_5_90_0)))))))) | (~i_2_5_99_0 & ((i_2_5_102_0 & ((i_2_5_62_0 & ((~i_2_5_65_0 & (i_2_5_12_0 | i_2_5_84_0 | ~i_2_5_90_0)) | (i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_90_0) | (i_2_5_12_0 & ((i_2_5_84_0 & ~i_2_5_90_0) | (i_2_5_82_0 & (i_2_5_84_0 | ~i_2_5_90_0)))))) | (~i_2_5_65_0 & ~i_2_5_90_0 & (i_2_5_12_0 | i_2_5_84_0)))) | (i_2_5_84_0 & ~i_2_5_90_0 & ((i_2_5_62_0 & ~i_2_5_65_0) | (i_2_5_12_0 & i_2_5_82_0))))) | (i_2_5_84_0 & ~i_2_5_90_0 & i_2_5_102_0 & i_2_5_12_0 & i_2_5_62_0 & ~i_2_5_65_0))) | (~i_2_5_90_0 & ((i_2_5_42_0 & ((i_2_5_12_0 & ((i_2_5_62_0 & ((~i_2_5_70_0 & (~i_2_5_91_0 | i_2_5_148_0)) | (~i_2_5_82_0 & ~i_2_5_84_0 & i_2_5_102_0 & ~i_2_5_148_0))) | (i_2_5_84_0 & ((~i_2_5_99_0 & i_2_5_102_0) | (i_2_5_82_0 & i_2_5_148_0))) | (~i_2_5_91_0 & ~i_2_5_99_0 & i_2_5_102_0) | (i_2_5_82_0 & ((~i_2_5_99_0 & i_2_5_102_0) | (~i_2_5_65_0 & ~i_2_5_84_0 & ~i_2_5_91_0))))) | (~i_2_5_65_0 & ((((i_2_5_84_0 & i_2_5_148_0) | (~i_2_5_70_0 & i_2_5_102_0)) & ((i_2_5_82_0 & ~i_2_5_91_0) | (i_2_5_62_0 & ~i_2_5_82_0))) | (i_2_5_82_0 & ((~i_2_5_70_0 & ((i_2_5_102_0 & i_2_5_148_0) | (i_2_5_84_0 & ~i_2_5_148_0))) | (i_2_5_84_0 & ((~i_2_5_91_0 & i_2_5_102_0) | (i_2_5_62_0 & ~i_2_5_102_0 & ~i_2_5_148_0))) | (~i_2_5_91_0 & ((i_2_5_62_0 & (i_2_5_102_0 | i_2_5_148_0)) | (i_2_5_102_0 & i_2_5_148_0))))) | (i_2_5_62_0 & ((~i_2_5_91_0 & ~i_2_5_99_0) | (~i_2_5_12_0 & ~i_2_5_70_0 & i_2_5_84_0))) | (~i_2_5_91_0 & ~i_2_5_99_0 & i_2_5_102_0) | (~i_2_5_70_0 & ((~i_2_5_91_0 & ~i_2_5_99_0) | (i_2_5_84_0 & i_2_5_102_0))))) | (i_2_5_62_0 & ((~i_2_5_70_0 & ((~i_2_5_91_0 & ~i_2_5_99_0) | (i_2_5_82_0 & i_2_5_84_0 & i_2_5_98_0 & ~i_2_5_102_0 & ~i_2_5_148_0))) | (i_2_5_82_0 & ((~i_2_5_99_0 & (i_2_5_148_0 | (i_2_5_84_0 & i_2_5_102_0))) | (~i_2_5_91_0 & ((i_2_5_102_0 & i_2_5_148_0) | (i_2_5_84_0 & (i_2_5_102_0 | i_2_5_148_0)))))) | (~i_2_5_91_0 & ((i_2_5_84_0 & (~i_2_5_99_0 | (i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_99_0 & (i_2_5_102_0 | i_2_5_148_0)))))) | (~i_2_5_91_0 & ((i_2_5_82_0 & ((i_2_5_84_0 & ((i_2_5_102_0 & i_2_5_148_0) | (~i_2_5_70_0 & (i_2_5_102_0 | i_2_5_148_0)))) | (~i_2_5_70_0 & ~i_2_5_99_0))) | (~i_2_5_99_0 & i_2_5_102_0 & (~i_2_5_70_0 | i_2_5_84_0 | i_2_5_148_0)))) | (~i_2_5_99_0 & i_2_5_102_0 & ~i_2_5_70_0 & i_2_5_82_0))) | ((~i_2_5_91_0 | (i_2_5_84_0 & i_2_5_102_0)) & ((i_2_5_12_0 & i_2_5_82_0 & ~i_2_5_99_0) | (i_2_5_62_0 & ~i_2_5_70_0 & i_2_5_148_0 & (~i_2_5_65_0 | i_2_5_82_0)))) | ((~i_2_5_70_0 | ~i_2_5_91_0) & ((~i_2_5_65_0 & ((i_2_5_12_0 & (~i_2_5_99_0 | (i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_99_0 & i_2_5_148_0) | (i_2_5_62_0 & i_2_5_102_0 & (~i_2_5_99_0 | (i_2_5_82_0 & i_2_5_84_0))))) | (i_2_5_84_0 & ((~i_2_5_99_0 & (i_2_5_12_0 | i_2_5_82_0)) | (i_2_5_12_0 & i_2_5_82_0 & (i_2_5_102_0 | i_2_5_148_0)))) | (i_2_5_102_0 & i_2_5_148_0 & i_2_5_12_0 & i_2_5_82_0))) | (~i_2_5_70_0 & ((i_2_5_12_0 & ((i_2_5_82_0 & ((i_2_5_84_0 & ~i_2_5_91_0) | (i_2_5_62_0 & ~i_2_5_65_0))) | ((~i_2_5_91_0 | i_2_5_102_0) & ((i_2_5_84_0 & i_2_5_148_0) | (i_2_5_62_0 & ~i_2_5_65_0))) | (~i_2_5_99_0 & i_2_5_102_0) | (~i_2_5_91_0 & ((i_2_5_102_0 & i_2_5_148_0) | ((i_2_5_62_0 | ~i_2_5_65_0) & (i_2_5_102_0 | i_2_5_148_0)))))) | (~i_2_5_99_0 & ((i_2_5_82_0 & (~i_2_5_65_0 | (~i_2_5_91_0 & i_2_5_102_0))) | (i_2_5_62_0 & ((~i_2_5_65_0 & (i_2_5_84_0 | ~i_2_5_91_0)) | (~i_2_5_91_0 & (i_2_5_84_0 | i_2_5_102_0)))) | (i_2_5_84_0 & i_2_5_102_0) | (~i_2_5_91_0 & (i_2_5_148_0 | (~i_2_5_65_0 & i_2_5_102_0))))) | (~i_2_5_91_0 & (((~i_2_5_65_0 | i_2_5_102_0) & ((i_2_5_82_0 & i_2_5_148_0) | (i_2_5_84_0 & (i_2_5_62_0 | i_2_5_148_0)))) | (i_2_5_102_0 & ((i_2_5_62_0 & (~i_2_5_65_0 | i_2_5_148_0)) | (~i_2_5_65_0 & i_2_5_148_0))) | (i_2_5_62_0 & i_2_5_84_0 & i_2_5_148_0))) | (~i_2_5_65_0 & i_2_5_82_0 & i_2_5_148_0 & ((i_2_5_62_0 & i_2_5_102_0) | (~i_2_5_42_0 & i_2_5_84_0))))) | (i_2_5_62_0 & ((~i_2_5_91_0 & (((i_2_5_84_0 | i_2_5_102_0) & ((~i_2_5_99_0 & i_2_5_148_0) | (~i_2_5_65_0 & (i_2_5_148_0 | (i_2_5_12_0 & i_2_5_82_0))))) | (i_2_5_12_0 & ((i_2_5_102_0 & i_2_5_148_0) | (~i_2_5_65_0 & (i_2_5_148_0 | (i_2_5_84_0 & i_2_5_102_0))))) | (i_2_5_102_0 & ((i_2_5_84_0 & ~i_2_5_99_0) | (i_2_5_82_0 & (~i_2_5_99_0 | (i_2_5_84_0 & i_2_5_148_0))))))) | (i_2_5_148_0 & ((i_2_5_12_0 & ((~i_2_5_65_0 & i_2_5_84_0) | (~i_2_5_82_0 & ~i_2_5_99_0))) | (~i_2_5_65_0 & i_2_5_82_0 & i_2_5_84_0 & i_2_5_102_0))) | (~i_2_5_65_0 & i_2_5_84_0 & ~i_2_5_99_0 & i_2_5_102_0))) | (i_2_5_84_0 & ((~i_2_5_65_0 & ~i_2_5_91_0 & (~i_2_5_99_0 | (i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_99_0 & i_2_5_148_0 & (i_2_5_12_0 | i_2_5_102_0)))) | (~i_2_5_99_0 & i_2_5_148_0 & i_2_5_82_0 & ~i_2_5_91_0))) | ((~i_2_5_91_0 | ~i_2_5_99_0) & ((i_2_5_148_0 & ((i_2_5_82_0 & ((i_2_5_62_0 & ~i_2_5_65_0 & ~i_2_5_70_0) | (i_2_5_12_0 & i_2_5_84_0 & i_2_5_102_0))) | (i_2_5_62_0 & ~i_2_5_65_0 & ~i_2_5_70_0 & (i_2_5_84_0 | i_2_5_102_0)))) | (~i_2_5_65_0 & ~i_2_5_70_0 & i_2_5_84_0 & i_2_5_102_0 & (i_2_5_62_0 | (~i_2_5_42_0 & ~i_2_5_82_0))))) | ((~i_2_5_99_0 | (~i_2_5_91_0 & i_2_5_102_0)) & ((i_2_5_12_0 & ~i_2_5_65_0 & ((i_2_5_62_0 & i_2_5_148_0) | (i_2_5_42_0 & i_2_5_84_0))) | (i_2_5_42_0 & i_2_5_62_0 & ~i_2_5_70_0 & i_2_5_82_0 & i_2_5_84_0))) | ((~i_2_5_91_0 | (i_2_5_62_0 & i_2_5_102_0)) & ((i_2_5_82_0 & ((i_2_5_12_0 & ~i_2_5_65_0 & i_2_5_84_0 & (~i_2_5_70_0 | i_2_5_148_0)) | (~i_2_5_70_0 & ~i_2_5_99_0 & i_2_5_148_0))) | (~i_2_5_65_0 & ~i_2_5_99_0 & i_2_5_12_0 & i_2_5_42_0))) | (~i_2_5_70_0 & (((~i_2_5_99_0 | i_2_5_148_0) & ((i_2_5_62_0 & ((i_2_5_12_0 & ((i_2_5_42_0 & i_2_5_84_0) | (~i_2_5_91_0 & i_2_5_102_0))) | (i_2_5_84_0 & ~i_2_5_91_0 & i_2_5_102_0))) | (i_2_5_84_0 & i_2_5_102_0 & i_2_5_12_0 & i_2_5_82_0))) | (i_2_5_62_0 & ((i_2_5_148_0 & ((i_2_5_12_0 & ((~i_2_5_65_0 & (~i_2_5_91_0 | (i_2_5_84_0 & i_2_5_102_0) | (i_2_5_82_0 & (i_2_5_84_0 | i_2_5_102_0)))) | (~i_2_5_99_0 & (i_2_5_84_0 | ~i_2_5_91_0)) | (i_2_5_42_0 & i_2_5_102_0))) | (~i_2_5_99_0 & ((~i_2_5_91_0 & i_2_5_102_0) | (i_2_5_42_0 & ~i_2_5_65_0))) | (i_2_5_82_0 & ((i_2_5_102_0 & ((~i_2_5_65_0 & i_2_5_84_0) | (i_2_5_42_0 & (~i_2_5_65_0 | ~i_2_5_91_0)))) | (i_2_5_42_0 & i_2_5_84_0 & ~i_2_5_91_0))) | (i_2_5_84_0 & i_2_5_102_0 & i_2_5_42_0 & ~i_2_5_82_0))) | (~i_2_5_91_0 & ((i_2_5_84_0 & ((~i_2_5_65_0 & ~i_2_5_99_0) | (i_2_5_12_0 & i_2_5_82_0 & i_2_5_102_0))) | (~i_2_5_65_0 & ((i_2_5_42_0 & (~i_2_5_99_0 | (i_2_5_82_0 & i_2_5_102_0))) | (~i_2_5_99_0 & (i_2_5_82_0 | i_2_5_102_0)))) | (~i_2_5_99_0 & i_2_5_102_0 & (i_2_5_42_0 | i_2_5_82_0)))) | (~i_2_5_99_0 & ((i_2_5_12_0 & ((~i_2_5_65_0 & i_2_5_102_0) | (i_2_5_42_0 & i_2_5_82_0))) | (~i_2_5_65_0 & i_2_5_82_0 & i_2_5_102_0))))) | (i_2_5_12_0 & ((~i_2_5_65_0 & ((i_2_5_84_0 & ~i_2_5_99_0) | (~i_2_5_91_0 & i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_91_0 & ((i_2_5_84_0 & ~i_2_5_99_0) | (i_2_5_82_0 & (~i_2_5_99_0 | (i_2_5_84_0 & i_2_5_148_0))) | (i_2_5_42_0 & (i_2_5_82_0 | (~i_2_5_99_0 & i_2_5_102_0))))) | (~i_2_5_99_0 & i_2_5_102_0 & (i_2_5_148_0 | (i_2_5_42_0 & i_2_5_82_0))))) | (i_2_5_84_0 & ((i_2_5_148_0 & (i_2_5_102_0 | (~i_2_5_65_0 & i_2_5_82_0)) & (~i_2_5_99_0 | (i_2_5_42_0 & ~i_2_5_91_0))) | (~i_2_5_99_0 & ((i_2_5_82_0 & ~i_2_5_91_0) | (i_2_5_42_0 & (~i_2_5_91_0 | (i_2_5_82_0 & i_2_5_102_0))))))) | (~i_2_5_65_0 & ~i_2_5_91_0 & ((i_2_5_82_0 & i_2_5_102_0 & i_2_5_148_0) | (~i_2_5_99_0 & (i_2_5_148_0 | (i_2_5_42_0 & (i_2_5_82_0 | i_2_5_102_0)))))) | (i_2_5_42_0 & i_2_5_90_0 & ~i_2_5_99_0 & i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_99_0 & ((i_2_5_12_0 & ((i_2_5_82_0 & ((i_2_5_42_0 & ((i_2_5_84_0 & ~i_2_5_91_0) | (i_2_5_102_0 & i_2_5_148_0))) | (i_2_5_62_0 & ((~i_2_5_65_0 & i_2_5_84_0) | (~i_2_5_91_0 & (i_2_5_102_0 | i_2_5_148_0)))))) | (~i_2_5_91_0 & ((i_2_5_102_0 & i_2_5_148_0) | (i_2_5_84_0 & (i_2_5_102_0 | i_2_5_148_0)) | (~i_2_5_65_0 & (i_2_5_62_0 | i_2_5_102_0)))) | (~i_2_5_65_0 & i_2_5_148_0 & (i_2_5_70_0 | i_2_5_102_0)))) | (~i_2_5_65_0 & (((i_2_5_84_0 | i_2_5_102_0) & ((~i_2_5_91_0 & i_2_5_148_0) | (i_2_5_62_0 & ((i_2_5_42_0 & ~i_2_5_91_0) | (i_2_5_82_0 & i_2_5_148_0))))) | (i_2_5_102_0 & ((i_2_5_84_0 & (~i_2_5_91_0 | i_2_5_148_0)) | (~i_2_5_42_0 & i_2_5_82_0 & ~i_2_5_91_0))))) | (~i_2_5_91_0 & ((i_2_5_148_0 & ((i_2_5_84_0 & i_2_5_102_0) | ((i_2_5_42_0 | i_2_5_82_0) & (i_2_5_84_0 | (i_2_5_62_0 & i_2_5_102_0))))) | (i_2_5_82_0 & i_2_5_84_0 & i_2_5_102_0))) | (i_2_5_42_0 & i_2_5_82_0 & i_2_5_84_0 & i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_91_0 & i_2_5_102_0 & ((i_2_5_148_0 & ((i_2_5_42_0 & ((i_2_5_12_0 & (i_2_5_62_0 | i_2_5_84_0)) | (i_2_5_62_0 & i_2_5_82_0 & (~i_2_5_65_0 | i_2_5_84_0)))) | (~i_2_5_65_0 & ((i_2_5_62_0 & i_2_5_84_0) | (i_2_5_12_0 & i_2_5_82_0))))) | (~i_2_5_65_0 & i_2_5_82_0 & i_2_5_84_0 & (i_2_5_12_0 | (i_2_5_42_0 & i_2_5_62_0))))))) | (~i_2_5_70_0 & ((i_2_5_62_0 & ((~i_2_5_90_0 & ((~i_2_5_12_0 & ((~i_2_5_84_0 & ~i_2_5_91_0 & ~i_2_5_98_0 & i_2_5_102_0) | (i_2_5_82_0 & i_2_5_84_0 & i_2_5_98_0 & ~i_2_5_99_0 & ~i_2_5_102_0))) | (i_2_5_82_0 & ((~i_2_5_84_0 & ~i_2_5_102_0 & ((i_2_5_12_0 & i_2_5_93_0 & ~i_2_5_99_0) | (i_2_5_42_0 & ~i_2_5_65_0 & i_2_5_148_0))) | ((i_2_5_102_0 | i_2_5_148_0) & ((i_2_5_12_0 & i_2_5_84_0 & ~i_2_5_91_0) | (~i_2_5_65_0 & ~i_2_5_98_0))) | (i_2_5_12_0 & ((~i_2_5_91_0 & i_2_5_102_0 & i_2_5_148_0) | (~i_2_5_98_0 & ~i_2_5_99_0))) | (i_2_5_84_0 & ((~i_2_5_98_0 & ((~i_2_5_91_0 & i_2_5_148_0) | (~i_2_5_99_0 & i_2_5_102_0))) | (~i_2_5_91_0 & (~i_2_5_65_0 | i_2_5_148_0) & (i_2_5_42_0 | i_2_5_102_0)) | (~i_2_5_65_0 & i_2_5_102_0 & i_2_5_148_0) | (i_2_5_42_0 & ~i_2_5_99_0))) | (i_2_5_102_0 & ((~i_2_5_98_0 & (~i_2_5_91_0 | i_2_5_148_0)) | (~i_2_5_91_0 & (~i_2_5_99_0 | (i_2_5_42_0 & i_2_5_148_0))))))) | ((i_2_5_12_0 | i_2_5_84_0) & ((~i_2_5_99_0 & i_2_5_148_0) | (~i_2_5_91_0 & ((~i_2_5_65_0 & i_2_5_148_0) | (~i_2_5_98_0 & ~i_2_5_99_0))))) | (~i_2_5_91_0 & (((~i_2_5_98_0 | i_2_5_102_0) & ((i_2_5_84_0 & ((i_2_5_42_0 & i_2_5_148_0) | (i_2_5_12_0 & ~i_2_5_65_0))) | (~i_2_5_65_0 & (~i_2_5_99_0 | i_2_5_148_0)))) | (~i_2_5_65_0 & ((i_2_5_42_0 & (~i_2_5_99_0 | (i_2_5_84_0 & i_2_5_102_0))) | (~i_2_5_98_0 & i_2_5_102_0) | (~i_2_5_99_0 & (i_2_5_84_0 | i_2_5_148_0)))) | (i_2_5_102_0 & ((i_2_5_84_0 & (~i_2_5_99_0 | (i_2_5_12_0 & i_2_5_148_0))) | (i_2_5_148_0 & (~i_2_5_98_0 | ~i_2_5_99_0)))) | (i_2_5_42_0 & ~i_2_5_98_0 & ~i_2_5_99_0))) | (~i_2_5_98_0 & ((i_2_5_148_0 & ((i_2_5_12_0 & (i_2_5_84_0 | i_2_5_102_0)) | ~i_2_5_99_0 | (~i_2_5_65_0 & i_2_5_102_0))) | (~i_2_5_65_0 & (i_2_5_42_0 | (i_2_5_84_0 & ~i_2_5_99_0))))) | (i_2_5_42_0 & i_2_5_102_0 & ((~i_2_5_82_0 & i_2_5_93_0 & ~i_2_5_99_0) | (~i_2_5_65_0 & i_2_5_84_0 & i_2_5_148_0))))) | (~i_2_5_98_0 & ((~i_2_5_148_0 & ((~i_2_5_65_0 & i_2_5_82_0 & ~i_2_5_84_0 & ~i_2_5_91_0 & i_2_5_93_0) | (i_2_5_12_0 & i_2_5_42_0 & i_2_5_91_0 & i_2_5_102_0))) | (~i_2_5_99_0 & (((~i_2_5_91_0 | i_2_5_102_0) & ((i_2_5_148_0 & (~i_2_5_65_0 | i_2_5_84_0)) | (~i_2_5_65_0 & (i_2_5_12_0 | i_2_5_42_0)))) | (((~i_2_5_91_0 & i_2_5_102_0) | (i_2_5_84_0 & (i_2_5_148_0 | (i_2_5_82_0 & i_2_5_102_0)))) & (i_2_5_42_0 | ~i_2_5_65_0)) | (i_2_5_12_0 & ((~i_2_5_65_0 & (i_2_5_148_0 | (i_2_5_82_0 & i_2_5_84_0))) | (~i_2_5_91_0 & (i_2_5_84_0 | i_2_5_102_0)) | (i_2_5_82_0 & (~i_2_5_91_0 | (i_2_5_84_0 & i_2_5_102_0))))) | (~i_2_5_91_0 & (((i_2_5_84_0 | i_2_5_148_0) & (i_2_5_82_0 | i_2_5_102_0)) | (i_2_5_82_0 & i_2_5_102_0) | (~i_2_5_65_0 & i_2_5_84_0))))) | (i_2_5_148_0 & ((~i_2_5_91_0 & (((i_2_5_82_0 | i_2_5_102_0) & (i_2_5_12_0 | i_2_5_42_0)) | (i_2_5_82_0 & i_2_5_84_0 & (~i_2_5_65_0 | i_2_5_102_0)))) | (~i_2_5_65_0 & i_2_5_82_0 & (i_2_5_42_0 | (i_2_5_84_0 & i_2_5_102_0))))) | (i_2_5_82_0 & ~i_2_5_91_0 & i_2_5_42_0 & ~i_2_5_65_0))) | (~i_2_5_91_0 & ((i_2_5_148_0 & (((i_2_5_82_0 | i_2_5_84_0) & ((~i_2_5_99_0 & i_2_5_102_0) | (i_2_5_12_0 & i_2_5_42_0))) | (i_2_5_102_0 & ((i_2_5_82_0 & ((i_2_5_42_0 & (~i_2_5_65_0 | i_2_5_84_0)) | (i_2_5_12_0 & i_2_5_84_0))) | (~i_2_5_65_0 & i_2_5_84_0) | (i_2_5_12_0 & (~i_2_5_65_0 | ~i_2_5_99_0)))) | (i_2_5_42_0 & (~i_2_5_99_0 | (~i_2_5_65_0 & i_2_5_82_0 & i_2_5_84_0))) | (~i_2_5_65_0 & i_2_5_84_0 & ~i_2_5_99_0))) | (i_2_5_82_0 & ((~i_2_5_65_0 & i_2_5_84_0 & ~i_2_5_99_0) | (i_2_5_102_0 & ((i_2_5_12_0 & (~i_2_5_65_0 | ~i_2_5_99_0)) | (i_2_5_84_0 & ~i_2_5_99_0) | (~i_2_5_65_0 & (~i_2_5_99_0 | (i_2_5_42_0 & i_2_5_84_0))))))) | (i_2_5_42_0 & ~i_2_5_99_0 & ((~i_2_5_65_0 & i_2_5_102_0) | (i_2_5_98_0 & ~i_2_5_102_0 & i_2_5_84_0 & i_2_5_90_0))))) | (~i_2_5_99_0 & ((i_2_5_12_0 & (i_2_5_42_0 | (i_2_5_84_0 & i_2_5_102_0)) & (i_2_5_148_0 | (~i_2_5_65_0 & i_2_5_82_0))) | (i_2_5_148_0 & ((i_2_5_42_0 & ((~i_2_5_65_0 & i_2_5_82_0) | (i_2_5_65_0 & i_2_5_102_0))) | (~i_2_5_65_0 & i_2_5_84_0 & i_2_5_102_0))))) | (i_2_5_84_0 & i_2_5_102_0 & i_2_5_148_0 & i_2_5_12_0 & i_2_5_42_0 & i_2_5_82_0))) | (~i_2_5_91_0 & (((~i_2_5_99_0 | (i_2_5_42_0 & i_2_5_148_0)) & ((i_2_5_82_0 & ((i_2_5_102_0 & ((i_2_5_12_0 & (~i_2_5_65_0 | ~i_2_5_90_0)) | (i_2_5_84_0 & (~i_2_5_90_0 | ~i_2_5_98_0)))) | (i_2_5_84_0 & ~i_2_5_90_0 & ~i_2_5_98_0))) | (i_2_5_12_0 & i_2_5_102_0 & ((~i_2_5_82_0 & i_2_5_84_0) | (~i_2_5_90_0 & ~i_2_5_98_0))))) | (~i_2_5_65_0 & ((~i_2_5_98_0 & ((i_2_5_93_0 & ~i_2_5_148_0 & ((~i_2_5_42_0 & i_2_5_82_0 & i_2_5_90_0 & i_2_5_102_0) | (i_2_5_12_0 & i_2_5_42_0 & ~i_2_5_102_0))) | ((i_2_5_82_0 | ~i_2_5_99_0) & ((i_2_5_42_0 & i_2_5_148_0) | (i_2_5_12_0 & i_2_5_102_0))) | ((~i_2_5_90_0 | i_2_5_102_0) & ((i_2_5_42_0 & ~i_2_5_99_0) | (i_2_5_148_0 & (i_2_5_12_0 | i_2_5_84_0)))) | (~i_2_5_90_0 & ((i_2_5_84_0 & ~i_2_5_99_0) | (i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_99_0 & ((i_2_5_102_0 & i_2_5_148_0) | (i_2_5_84_0 & (i_2_5_42_0 | i_2_5_148_0)))))) | (i_2_5_42_0 & ((~i_2_5_90_0 & (((i_2_5_102_0 | i_2_5_148_0) & (~i_2_5_99_0 | (i_2_5_12_0 & i_2_5_82_0))) | (i_2_5_84_0 & ~i_2_5_99_0) | (i_2_5_148_0 & ((i_2_5_82_0 & (i_2_5_84_0 | i_2_5_102_0)) | (i_2_5_12_0 & i_2_5_84_0))))) | (i_2_5_148_0 & ((~i_2_5_99_0 & i_2_5_102_0) | (i_2_5_84_0 & (~i_2_5_99_0 | (i_2_5_82_0 & i_2_5_102_0))))) | (i_2_5_12_0 & ~i_2_5_99_0 & i_2_5_102_0))) | (i_2_5_12_0 & ((i_2_5_82_0 & i_2_5_84_0 & (~i_2_5_90_0 | i_2_5_148_0)) | (~i_2_5_99_0 & i_2_5_102_0 & i_2_5_148_0) | (~i_2_5_90_0 & (~i_2_5_99_0 | (i_2_5_102_0 & i_2_5_148_0))))) | (i_2_5_84_0 & i_2_5_102_0 & (~i_2_5_99_0 | (~i_2_5_90_0 & i_2_5_148_0))))) | (~i_2_5_98_0 & ((~i_2_5_90_0 & ((i_2_5_82_0 & ((~i_2_5_42_0 & (~i_2_5_99_0 | (i_2_5_84_0 & i_2_5_102_0))) | (i_2_5_42_0 & ~i_2_5_84_0 & i_2_5_102_0))) | (~i_2_5_99_0 & ((i_2_5_102_0 & i_2_5_148_0) | ((i_2_5_102_0 | i_2_5_148_0) & (i_2_5_42_0 | i_2_5_84_0)))))) | (~i_2_5_99_0 & ((i_2_5_102_0 & ((i_2_5_12_0 & (i_2_5_82_0 | i_2_5_148_0)) | (i_2_5_148_0 & (i_2_5_42_0 | i_2_5_84_0)))) | (i_2_5_42_0 & i_2_5_84_0 & i_2_5_148_0))) | (i_2_5_12_0 & i_2_5_82_0 & ((i_2_5_84_0 & i_2_5_102_0) | (i_2_5_42_0 & i_2_5_148_0))))) | (i_2_5_148_0 & ((i_2_5_12_0 & ((i_2_5_82_0 & (~i_2_5_99_0 | (i_2_5_84_0 & ~i_2_5_90_0 & i_2_5_102_0))) | (~i_2_5_99_0 & (i_2_5_42_0 | i_2_5_84_0)))) | (~i_2_5_99_0 & ((i_2_5_82_0 & i_2_5_84_0) | (i_2_5_42_0 & ((~i_2_5_90_0 & i_2_5_102_0) | (i_2_5_84_0 & (~i_2_5_90_0 | i_2_5_102_0)))))))) | (i_2_5_12_0 & ~i_2_5_90_0 & ~i_2_5_99_0 & (i_2_5_42_0 | i_2_5_84_0)))) | (i_2_5_102_0 & ((i_2_5_84_0 & ((i_2_5_42_0 & ((i_2_5_82_0 & ((i_2_5_12_0 & (~i_2_5_99_0 | (~i_2_5_90_0 & i_2_5_148_0))) | (~i_2_5_99_0 & i_2_5_148_0) | (~i_2_5_65_0 & ~i_2_5_90_0 & ~i_2_5_148_0))) | (~i_2_5_65_0 & ((~i_2_5_98_0 & ~i_2_5_99_0) | (i_2_5_12_0 & ~i_2_5_90_0 & ~i_2_5_148_0))) | (~i_2_5_90_0 & ~i_2_5_98_0 & (~i_2_5_82_0 | ~i_2_5_99_0)))) | (~i_2_5_99_0 & ((i_2_5_12_0 & (~i_2_5_90_0 | (~i_2_5_65_0 & i_2_5_82_0 & ~i_2_5_98_0))) | (i_2_5_148_0 & (~i_2_5_90_0 | (~i_2_5_42_0 & ~i_2_5_65_0 & ~i_2_5_82_0))))) | (~i_2_5_90_0 & ~i_2_5_98_0 & i_2_5_12_0 & ~i_2_5_82_0))) | (~i_2_5_99_0 & ((i_2_5_12_0 & ((i_2_5_42_0 & i_2_5_82_0 & (i_2_5_148_0 | (~i_2_5_65_0 & ~i_2_5_98_0))) | (i_2_5_148_0 & (~i_2_5_90_0 | (~i_2_5_65_0 & ~i_2_5_98_0))))) | (~i_2_5_65_0 & ((~i_2_5_90_0 & ~i_2_5_98_0) | (i_2_5_82_0 & (~i_2_5_90_0 | (i_2_5_42_0 & ~i_2_5_98_0 & i_2_5_148_0))))))) | (~i_2_5_90_0 & ~i_2_5_98_0 & ((i_2_5_42_0 & ~i_2_5_65_0) | (i_2_5_12_0 & i_2_5_82_0 & i_2_5_148_0))))) | (~i_2_5_98_0 & ((i_2_5_82_0 & ((~i_2_5_90_0 & ((i_2_5_12_0 & i_2_5_84_0 & ~i_2_5_102_0) | (i_2_5_42_0 & ~i_2_5_65_0 & ~i_2_5_148_0))) | (~i_2_5_99_0 & ((i_2_5_148_0 & ((~i_2_5_65_0 & i_2_5_84_0) | (i_2_5_12_0 & (i_2_5_42_0 | i_2_5_84_0)))) | (i_2_5_42_0 & ~i_2_5_65_0 & i_2_5_84_0))))) | (i_2_5_12_0 & i_2_5_42_0 & i_2_5_65_0 & i_2_5_84_0 & ~i_2_5_90_0))) | (i_2_5_12_0 & ~i_2_5_90_0 & i_2_5_91_0 & ~i_2_5_99_0 & i_2_5_148_0))) | (~i_2_5_98_0 & ((i_2_5_62_0 & ((~i_2_5_65_0 & ((~i_2_5_12_0 & ((i_2_5_70_0 & i_2_5_82_0 & ~i_2_5_84_0 & ~i_2_5_99_0 & ~i_2_5_102_0 & i_2_5_148_0) | (i_2_5_42_0 & i_2_5_84_0 & ~i_2_5_90_0 & i_2_5_93_0 & ~i_2_5_148_0))) | (i_2_5_148_0 & ((~i_2_5_82_0 & ((i_2_5_12_0 & i_2_5_84_0 & i_2_5_102_0) | (i_2_5_42_0 & ~i_2_5_91_0 & i_2_5_93_0))) | (i_2_5_12_0 & ((i_2_5_84_0 & ~i_2_5_91_0) | (i_2_5_82_0 & ~i_2_5_84_0 & i_2_5_102_0))) | (i_2_5_42_0 & ((~i_2_5_99_0 & i_2_5_102_0) | (i_2_5_84_0 & ~i_2_5_90_0 & ~i_2_5_102_0))) | (~i_2_5_90_0 & (~i_2_5_99_0 | (~i_2_5_91_0 & i_2_5_102_0))) | (~i_2_5_91_0 & ((i_2_5_84_0 & ~i_2_5_99_0) | (~i_2_5_84_0 & i_2_5_102_0))))) | (i_2_5_93_0 & ((i_2_5_42_0 & ~i_2_5_90_0 & ~i_2_5_99_0) | (~i_2_5_91_0 & i_2_5_102_0 & i_2_5_82_0 & i_2_5_90_0))) | (~i_2_5_99_0 & ((i_2_5_84_0 & ((i_2_5_12_0 & (i_2_5_42_0 | (i_2_5_82_0 & i_2_5_102_0))) | (~i_2_5_91_0 & (~i_2_5_90_0 | i_2_5_102_0)) | (i_2_5_42_0 & i_2_5_82_0 & ~i_2_5_102_0))) | (~i_2_5_90_0 & ((~i_2_5_91_0 & i_2_5_102_0) | (i_2_5_12_0 & ~i_2_5_102_0))) | (i_2_5_42_0 & ~i_2_5_91_0 & i_2_5_102_0))) | (~i_2_5_91_0 & ((i_2_5_102_0 & ((i_2_5_12_0 & i_2_5_82_0) | ((i_2_5_42_0 | i_2_5_84_0) & (i_2_5_12_0 | i_2_5_82_0)))) | (i_2_5_42_0 & i_2_5_84_0 & ~i_2_5_90_0))) | (i_2_5_82_0 & ~i_2_5_90_0 & ((i_2_5_84_0 & i_2_5_102_0) | (i_2_5_12_0 & ~i_2_5_84_0))))) | (i_2_5_102_0 & ((i_2_5_84_0 & ((i_2_5_12_0 & ((~i_2_5_82_0 & ((~i_2_5_90_0 & i_2_5_148_0) | (i_2_5_42_0 & i_2_5_90_0 & ~i_2_5_91_0))) | (~i_2_5_91_0 & (~i_2_5_99_0 | (i_2_5_82_0 & i_2_5_148_0))) | (i_2_5_82_0 & ~i_2_5_99_0 & (~i_2_5_90_0 | i_2_5_148_0)))) | (~i_2_5_91_0 & ((i_2_5_42_0 & ((i_2_5_82_0 & ~i_2_5_99_0) | (~i_2_5_90_0 & i_2_5_148_0))) | (~i_2_5_99_0 & i_2_5_148_0) | (~i_2_5_90_0 & (~i_2_5_99_0 | (i_2_5_82_0 & i_2_5_148_0))))) | (i_2_5_42_0 & ~i_2_5_99_0 & (i_2_5_148_0 | (~i_2_5_82_0 & ~i_2_5_90_0))))) | (~i_2_5_91_0 & ((i_2_5_82_0 & ((~i_2_5_99_0 & (~i_2_5_90_0 | i_2_5_148_0)) | (i_2_5_42_0 & ((i_2_5_12_0 & ~i_2_5_99_0) | (~i_2_5_90_0 & i_2_5_148_0))))) | (~i_2_5_99_0 & i_2_5_148_0 & (i_2_5_42_0 | ~i_2_5_90_0)))))) | (~i_2_5_91_0 & ((~i_2_5_99_0 & ((i_2_5_12_0 & (i_2_5_148_0 | (i_2_5_84_0 & ~i_2_5_90_0))) | (~i_2_5_90_0 & ((i_2_5_84_0 & i_2_5_148_0) | (i_2_5_42_0 & (i_2_5_148_0 | (i_2_5_82_0 & i_2_5_84_0))))) | (i_2_5_82_0 & i_2_5_84_0 & i_2_5_148_0))) | (i_2_5_12_0 & ~i_2_5_42_0 & i_2_5_82_0 & ~i_2_5_90_0 & i_2_5_148_0))) | (~i_2_5_99_0 & i_2_5_148_0 & i_2_5_12_0 & ~i_2_5_90_0))) | (~i_2_5_99_0 & ((~i_2_5_65_0 & ((i_2_5_84_0 & ((~i_2_5_91_0 & ((i_2_5_12_0 & (~i_2_5_42_0 | ~i_2_5_90_0)) | i_2_5_82_0 | (~i_2_5_90_0 & i_2_5_102_0))) | (i_2_5_148_0 & ((i_2_5_42_0 & (i_2_5_82_0 | i_2_5_102_0)) | (i_2_5_82_0 & i_2_5_102_0) | (~i_2_5_42_0 & ~i_2_5_90_0))))) | (i_2_5_12_0 & ((i_2_5_82_0 & (~i_2_5_91_0 | (i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_91_0 & (i_2_5_148_0 | (~i_2_5_90_0 & i_2_5_102_0))))) | (i_2_5_42_0 & ~i_2_5_91_0 & ((i_2_5_102_0 & i_2_5_148_0) | (~i_2_5_90_0 & (i_2_5_102_0 | i_2_5_148_0)))) | (~i_2_5_90_0 & i_2_5_102_0 & i_2_5_148_0))) | (~i_2_5_91_0 & ((~i_2_5_90_0 & ((i_2_5_12_0 & ((i_2_5_82_0 & i_2_5_102_0) | (~i_2_5_42_0 & i_2_5_148_0))) | (i_2_5_82_0 & i_2_5_84_0 & i_2_5_148_0) | (i_2_5_102_0 & ((i_2_5_84_0 & i_2_5_148_0) | (i_2_5_42_0 & (i_2_5_148_0 | (i_2_5_82_0 & i_2_5_84_0))))))) | (i_2_5_82_0 & i_2_5_148_0 & ((i_2_5_84_0 & i_2_5_102_0) | (i_2_5_12_0 & (~i_2_5_42_0 | i_2_5_102_0)))))) | (i_2_5_82_0 & ~i_2_5_90_0 & i_2_5_102_0 & i_2_5_148_0 & (i_2_5_42_0 | i_2_5_84_0)))) | (~i_2_5_91_0 & ((~i_2_5_90_0 & ((i_2_5_82_0 & ((i_2_5_42_0 & ((~i_2_5_65_0 & i_2_5_102_0) | (i_2_5_12_0 & i_2_5_84_0 & ~i_2_5_148_0))) | (i_2_5_12_0 & (~i_2_5_65_0 | (i_2_5_84_0 & i_2_5_102_0))) | (~i_2_5_65_0 & ((i_2_5_84_0 & i_2_5_102_0) | (~i_2_5_102_0 & i_2_5_148_0))))) | (i_2_5_102_0 & i_2_5_148_0 & ((i_2_5_42_0 & ~i_2_5_65_0 & i_2_5_84_0) | (i_2_5_12_0 & ((~i_2_5_65_0 & i_2_5_84_0) | (i_2_5_42_0 & (~i_2_5_65_0 | i_2_5_84_0)))))))) | (i_2_5_12_0 & ~i_2_5_65_0 & ((i_2_5_82_0 & (i_2_5_84_0 | (i_2_5_70_0 & i_2_5_148_0))) | (i_2_5_42_0 & i_2_5_84_0 & i_2_5_102_0))))) | (i_2_5_12_0 & i_2_5_42_0 & i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_90_0 & i_2_5_99_0 & i_2_5_102_0))) | (~i_2_5_99_0 & ((~i_2_5_91_0 & (((i_2_5_84_0 | i_2_5_102_0) & ((i_2_5_12_0 & i_2_5_62_0 & ~i_2_5_65_0) | (~i_2_5_90_0 & i_2_5_148_0 & ~i_2_5_42_0 & i_2_5_82_0))) | (i_2_5_102_0 & (((i_2_5_62_0 | i_2_5_84_0) & ((~i_2_5_65_0 & i_2_5_148_0) | (i_2_5_12_0 & ~i_2_5_82_0 & ~i_2_5_90_0))) | (~i_2_5_65_0 & ((i_2_5_42_0 & ((i_2_5_12_0 & i_2_5_148_0) | (i_2_5_62_0 & ~i_2_5_90_0))) | (i_2_5_82_0 & (i_2_5_84_0 | i_2_5_148_0)) | (~i_2_5_90_0 & (i_2_5_148_0 | (i_2_5_62_0 & i_2_5_84_0))))) | (i_2_5_12_0 & ((i_2_5_42_0 & ((i_2_5_82_0 & i_2_5_84_0) | (i_2_5_62_0 & ~i_2_5_90_0))) | (i_2_5_84_0 & i_2_5_148_0) | (i_2_5_62_0 & ((i_2_5_84_0 & ~i_2_5_90_0) | (i_2_5_82_0 & i_2_5_148_0))))) | (i_2_5_84_0 & ((i_2_5_82_0 & ~i_2_5_90_0 & i_2_5_148_0) | (i_2_5_62_0 & ((~i_2_5_90_0 & i_2_5_148_0) | (i_2_5_82_0 & (i_2_5_148_0 | (i_2_5_42_0 & ~i_2_5_90_0))))))))) | (i_2_5_148_0 & ((~i_2_5_65_0 & ((i_2_5_12_0 & (i_2_5_62_0 | ~i_2_5_90_0)) | ((i_2_5_82_0 | (i_2_5_84_0 & ~i_2_5_90_0)) & (i_2_5_42_0 | i_2_5_62_0)))) | (i_2_5_12_0 & ~i_2_5_90_0 & (i_2_5_82_0 | i_2_5_84_0)))) | (i_2_5_62_0 & i_2_5_82_0 & ((~i_2_5_65_0 & ~i_2_5_90_0) | (i_2_5_12_0 & i_2_5_42_0 & i_2_5_84_0))))) | (~i_2_5_65_0 & ((i_2_5_62_0 & ((i_2_5_42_0 & ((i_2_5_82_0 & i_2_5_84_0 & i_2_5_98_0 & i_2_5_102_0) | (i_2_5_70_0 & ~i_2_5_90_0 & i_2_5_93_0 & i_2_5_148_0))) | (i_2_5_102_0 & i_2_5_148_0 & (~i_2_5_90_0 | (i_2_5_12_0 & i_2_5_98_0))))) | (~i_2_5_90_0 & ((i_2_5_82_0 & i_2_5_148_0) | (i_2_5_12_0 & (i_2_5_82_0 | (i_2_5_84_0 & i_2_5_102_0))))))) | (i_2_5_62_0 & ((i_2_5_12_0 & ((~i_2_5_90_0 & i_2_5_102_0 & i_2_5_148_0) | (i_2_5_42_0 & ~i_2_5_84_0 & ((i_2_5_102_0 & i_2_5_148_0) | (i_2_5_82_0 & ~i_2_5_90_0 & ~i_2_5_102_0))))) | (i_2_5_42_0 & ~i_2_5_90_0 & i_2_5_93_0 & i_2_5_98_0 & i_2_5_102_0 & i_2_5_148_0))))) | (~i_2_5_65_0 & ((~i_2_5_90_0 & ((i_2_5_42_0 & ((i_2_5_62_0 & ((i_2_5_12_0 & ((i_2_5_82_0 & i_2_5_148_0) | (~i_2_5_82_0 & ~i_2_5_91_0 & i_2_5_99_0))) | (~i_2_5_91_0 & i_2_5_148_0 & ((i_2_5_84_0 & i_2_5_102_0) | (i_2_5_82_0 & (i_2_5_84_0 | i_2_5_102_0)))))) | (~i_2_5_91_0 & i_2_5_102_0 & i_2_5_148_0 & ((i_2_5_82_0 & i_2_5_84_0) | (i_2_5_12_0 & (i_2_5_82_0 | i_2_5_84_0)))))) | (i_2_5_84_0 & ~i_2_5_91_0 & ((i_2_5_12_0 & ((i_2_5_62_0 & i_2_5_102_0 & (i_2_5_82_0 | i_2_5_148_0)) | (~i_2_5_42_0 & i_2_5_82_0 & i_2_5_148_0))) | (i_2_5_62_0 & i_2_5_82_0 & i_2_5_102_0 & i_2_5_148_0))))) | (i_2_5_12_0 & i_2_5_62_0 & ~i_2_5_91_0 & i_2_5_148_0 & ((i_2_5_42_0 & i_2_5_84_0 & i_2_5_102_0) | (i_2_5_82_0 & i_2_5_93_0))))) | (i_2_5_12_0 & i_2_5_62_0 & i_2_5_84_0 & ~i_2_5_90_0 & ~i_2_5_91_0 & i_2_5_102_0 & i_2_5_148_0 & (i_2_5_42_0 | i_2_5_82_0)))) | (~i_2_5_91_0 & ((~i_2_5_93_0 & ((i_2_5_102_0 & ((i_2_5_84_0 & ((~i_2_5_42_0 & ((i_2_5_62_0 & i_2_5_82_0 & ~i_2_5_90_0 & ~i_2_5_99_0) | (~i_2_5_65_0 & ~i_2_5_70_0 & i_2_5_148_0))) | (((i_2_5_12_0 & ~i_2_5_65_0) | (i_2_5_82_0 & ~i_2_5_98_0 & i_2_5_148_0)) & ((i_2_5_62_0 & ~i_2_5_99_0) | (~i_2_5_62_0 & ~i_2_5_70_0))) | (i_2_5_62_0 & ((~i_2_5_99_0 & (((~i_2_5_70_0 | ~i_2_5_90_0) & (i_2_5_12_0 | (~i_2_5_65_0 & ~i_2_5_98_0))) | (~i_2_5_65_0 & (i_2_5_82_0 | (i_2_5_42_0 & ~i_2_5_98_0))) | (i_2_5_148_0 & (~i_2_5_90_0 | (i_2_5_42_0 & ~i_2_5_98_0))) | (i_2_5_42_0 & ((~i_2_5_90_0 & ~i_2_5_98_0) | (~i_2_5_70_0 & ~i_2_5_82_0))) | (~i_2_5_70_0 & ~i_2_5_98_0 & (i_2_5_82_0 | ~i_2_5_90_0)))) | (~i_2_5_90_0 & ((i_2_5_42_0 & ((~i_2_5_70_0 & i_2_5_82_0) | (~i_2_5_98_0 & i_2_5_148_0) | (~i_2_5_65_0 & i_2_5_70_0 & ~i_2_5_82_0 & i_2_5_98_0 & ~i_2_5_148_0))) | (~i_2_5_98_0 & ((~i_2_5_70_0 & i_2_5_148_0) | (~i_2_5_65_0 & (~i_2_5_70_0 | i_2_5_148_0)))))))) | (~i_2_5_90_0 & ((i_2_5_42_0 & ((~i_2_5_82_0 & ((~i_2_5_70_0 & ~i_2_5_99_0) | (i_2_5_12_0 & ~i_2_5_98_0 & i_2_5_99_0))) | (~i_2_5_99_0 & (i_2_5_148_0 | (~i_2_5_65_0 & ~i_2_5_98_0))))) | (i_2_5_12_0 & ((~i_2_5_65_0 & (~i_2_5_99_0 | (i_2_5_82_0 & ~i_2_5_98_0))) | (i_2_5_82_0 & ~i_2_5_98_0 & i_2_5_148_0) | (~i_2_5_70_0 & (i_2_5_148_0 | (i_2_5_82_0 & ~i_2_5_98_0))))) | (i_2_5_82_0 & ~i_2_5_99_0 & (~i_2_5_65_0 | (~i_2_5_70_0 & ~i_2_5_98_0))))) | (i_2_5_82_0 & ((~i_2_5_65_0 & ((i_2_5_42_0 & ~i_2_5_70_0) | (i_2_5_90_0 & i_2_5_148_0))) | (i_2_5_12_0 & ~i_2_5_98_0 & ~i_2_5_99_0))) | (~i_2_5_70_0 & ((i_2_5_12_0 & (i_2_5_42_0 | (~i_2_5_98_0 & i_2_5_148_0))) | (i_2_5_42_0 & ~i_2_5_99_0 & i_2_5_148_0))) | (i_2_5_12_0 & ~i_2_5_99_0 & i_2_5_148_0))) | (~i_2_5_65_0 & ((~i_2_5_82_0 & ((i_2_5_62_0 & ~i_2_5_70_0 & ~i_2_5_84_0 & ~i_2_5_90_0 & i_2_5_98_0) | (i_2_5_12_0 & ~i_2_5_42_0 & i_2_5_90_0 & ~i_2_5_98_0 & i_2_5_148_0))) | (i_2_5_148_0 & ((~i_2_5_70_0 & ((~i_2_5_12_0 & ((i_2_5_42_0 & ~i_2_5_98_0) | (~i_2_5_42_0 & i_2_5_62_0 & i_2_5_98_0))) | (~i_2_5_90_0 & ~i_2_5_99_0) | (i_2_5_62_0 & (~i_2_5_90_0 | (i_2_5_12_0 & ~i_2_5_98_0))))) | (i_2_5_12_0 & ((~i_2_5_98_0 & ~i_2_5_99_0) | (i_2_5_62_0 & ~i_2_5_90_0))) | (i_2_5_62_0 & ~i_2_5_99_0) | (~i_2_5_98_0 & ((~i_2_5_90_0 & (i_2_5_82_0 | ~i_2_5_99_0)) | (~i_2_5_42_0 & ~i_2_5_99_0))))) | (i_2_5_42_0 & ((i_2_5_82_0 & ((i_2_5_12_0 & i_2_5_62_0) | (~i_2_5_12_0 & i_2_5_70_0 & ~i_2_5_84_0 & ~i_2_5_90_0 & ~i_2_5_98_0))) | (~i_2_5_99_0 & ((~i_2_5_98_0 & (~i_2_5_70_0 | ~i_2_5_90_0) & (i_2_5_12_0 | i_2_5_62_0)) | (i_2_5_12_0 & ~i_2_5_70_0 & ~i_2_5_90_0))))) | (i_2_5_62_0 & ((~i_2_5_70_0 & (((~i_2_5_90_0 | ~i_2_5_99_0) & (i_2_5_12_0 | (i_2_5_82_0 & ~i_2_5_98_0))) | (~i_2_5_90_0 & ~i_2_5_99_0) | (i_2_5_12_0 & i_2_5_98_0 & ~i_2_5_148_0))) | (~i_2_5_99_0 & ((i_2_5_12_0 & (i_2_5_82_0 | ~i_2_5_90_0)) | (i_2_5_82_0 & ~i_2_5_90_0))))) | (~i_2_5_70_0 & ~i_2_5_99_0 & ((i_2_5_12_0 & i_2_5_82_0) | (~i_2_5_90_0 & ~i_2_5_98_0))))) | (~i_2_5_70_0 & ((~i_2_5_90_0 & ((i_2_5_42_0 & ((i_2_5_62_0 & ((~i_2_5_12_0 & i_2_5_65_0 & ~i_2_5_84_0 & ~i_2_5_98_0) | (i_2_5_82_0 & ~i_2_5_148_0))) | (~i_2_5_99_0 & ((i_2_5_82_0 & ~i_2_5_84_0) | (i_2_5_12_0 & ~i_2_5_98_0))))) | (i_2_5_12_0 & ((i_2_5_62_0 & ~i_2_5_99_0) | (~i_2_5_98_0 & i_2_5_148_0))) | (~i_2_5_98_0 & ~i_2_5_99_0 & (i_2_5_148_0 | (i_2_5_62_0 & i_2_5_82_0))))) | (~i_2_5_99_0 & ((i_2_5_12_0 & (i_2_5_148_0 | (i_2_5_62_0 & i_2_5_82_0))) | (i_2_5_82_0 & (i_2_5_148_0 | (i_2_5_42_0 & i_2_5_62_0 & ~i_2_5_98_0))))))) | (~i_2_5_99_0 & ((i_2_5_62_0 & ((i_2_5_42_0 & ((i_2_5_12_0 & ~i_2_5_90_0) | (i_2_5_82_0 & ~i_2_5_98_0 & i_2_5_148_0))) | (i_2_5_12_0 & i_2_5_82_0 & (~i_2_5_90_0 | i_2_5_148_0)))) | (~i_2_5_90_0 & ~i_2_5_98_0 & i_2_5_148_0 & (i_2_5_12_0 | i_2_5_82_0)))))) | (~i_2_5_99_0 & ((~i_2_5_70_0 & ((i_2_5_62_0 & ((i_2_5_98_0 & ((i_2_5_12_0 & ~i_2_5_82_0 & ~i_2_5_90_0) | (~i_2_5_12_0 & ~i_2_5_102_0 & ((i_2_5_84_0 & i_2_5_148_0) | (i_2_5_65_0 & i_2_5_82_0 & ~i_2_5_84_0 & ~i_2_5_90_0))))) | (~i_2_5_98_0 & ((i_2_5_82_0 & ((i_2_5_84_0 & ~i_2_5_90_0) | (i_2_5_12_0 & ~i_2_5_65_0))) | (~i_2_5_65_0 & (~i_2_5_90_0 | i_2_5_148_0)) | (~i_2_5_90_0 & (i_2_5_148_0 | (i_2_5_42_0 & i_2_5_84_0))))) | (~i_2_5_65_0 & i_2_5_82_0 & i_2_5_84_0) | (~i_2_5_90_0 & ((i_2_5_42_0 & i_2_5_82_0) | (i_2_5_12_0 & (i_2_5_42_0 | i_2_5_84_0)))))) | (i_2_5_12_0 & ((i_2_5_42_0 & (i_2_5_84_0 | (~i_2_5_65_0 & ~i_2_5_90_0 & ~i_2_5_98_0))) | (~i_2_5_98_0 & ((i_2_5_82_0 & (i_2_5_84_0 | ~i_2_5_90_0)) | (i_2_5_84_0 & (~i_2_5_65_0 | i_2_5_148_0)))))) | (~i_2_5_98_0 & ((i_2_5_84_0 & ((i_2_5_42_0 & (~i_2_5_65_0 | i_2_5_148_0)) | (~i_2_5_65_0 & i_2_5_82_0 & ~i_2_5_90_0))) | (i_2_5_148_0 & (i_2_5_82_0 | (~i_2_5_65_0 & ~i_2_5_90_0))))) | (~i_2_5_65_0 & i_2_5_84_0 & ~i_2_5_90_0 & i_2_5_148_0))) | (~i_2_5_65_0 & ((~i_2_5_90_0 & ((i_2_5_42_0 & ~i_2_5_98_0 & (i_2_5_82_0 | (i_2_5_62_0 & i_2_5_84_0))) | (~i_2_5_42_0 & ((i_2_5_84_0 & i_2_5_148_0) | (i_2_5_12_0 & i_2_5_82_0))) | (i_2_5_62_0 & i_2_5_148_0) | ((i_2_5_12_0 | i_2_5_82_0) & (i_2_5_148_0 | (i_2_5_62_0 & i_2_5_84_0))))) | (i_2_5_12_0 & ((i_2_5_82_0 & i_2_5_84_0) | (i_2_5_62_0 & i_2_5_148_0))) | (i_2_5_148_0 & ((i_2_5_42_0 & ((i_2_5_62_0 & i_2_5_70_0 & ~i_2_5_84_0 & i_2_5_98_0) | (i_2_5_84_0 & ~i_2_5_98_0))) | (i_2_5_70_0 & i_2_5_82_0))) | (i_2_5_42_0 & i_2_5_82_0 & i_2_5_84_0))) | (~i_2_5_90_0 & ((i_2_5_84_0 & ((i_2_5_12_0 & (i_2_5_148_0 | (i_2_5_82_0 & ~i_2_5_98_0))) | (i_2_5_62_0 & i_2_5_148_0 & (i_2_5_42_0 | i_2_5_82_0)))) | (i_2_5_82_0 & i_2_5_148_0 & i_2_5_42_0 & i_2_5_62_0))) | (i_2_5_12_0 & i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_98_0 & i_2_5_148_0))) | (i_2_5_42_0 & ((i_2_5_82_0 & ((~i_2_5_98_0 & ((i_2_5_12_0 & i_2_5_90_0 & i_2_5_99_0 & ((i_2_5_62_0 & i_2_5_84_0) | (~i_2_5_65_0 & i_2_5_70_0))) | (i_2_5_62_0 & ~i_2_5_65_0 & ~i_2_5_90_0 & ~i_2_5_148_0))) | (i_2_5_62_0 & ~i_2_5_65_0 & ((~i_2_5_70_0 & (i_2_5_84_0 | (~i_2_5_90_0 & ~i_2_5_148_0))) | (i_2_5_84_0 & i_2_5_148_0 & (~i_2_5_90_0 | i_2_5_98_0)))))) | (i_2_5_84_0 & ((i_2_5_12_0 & i_2_5_148_0 & ((i_2_5_62_0 & ~i_2_5_90_0) | (~i_2_5_65_0 & i_2_5_90_0))) | (~i_2_5_90_0 & ~i_2_5_102_0 & ~i_2_5_148_0 & i_2_5_62_0 & ~i_2_5_65_0 & ~i_2_5_70_0))) | (i_2_5_62_0 & ~i_2_5_70_0 & ~i_2_5_84_0 & ~i_2_5_90_0 & ~i_2_5_98_0 & i_2_5_148_0))) | (~i_2_5_65_0 & ((~i_2_5_70_0 & ((i_2_5_84_0 & ((i_2_5_12_0 & ((~i_2_5_98_0 & i_2_5_148_0) | (i_2_5_62_0 & ~i_2_5_90_0))) | (~i_2_5_90_0 & i_2_5_148_0 & ((~i_2_5_42_0 & i_2_5_82_0) | (i_2_5_62_0 & ~i_2_5_98_0))))) | (~i_2_5_98_0 & i_2_5_148_0 & i_2_5_12_0 & ~i_2_5_90_0))) | (~i_2_5_90_0 & i_2_5_148_0 & i_2_5_12_0 & i_2_5_82_0))) | (~i_2_5_90_0 & ~i_2_5_98_0 & i_2_5_148_0 & i_2_5_12_0 & ~i_2_5_70_0 & i_2_5_84_0))) | (~i_2_5_70_0 & ((i_2_5_102_0 & ((i_2_5_148_0 & ((~i_2_5_42_0 & ((~i_2_5_65_0 & i_2_5_84_0 & i_2_5_12_0 & i_2_5_62_0) | (~i_2_5_98_0 & ~i_2_5_99_0 & i_2_5_82_0 & i_2_5_90_0))) | (i_2_5_62_0 & ((i_2_5_12_0 & ((~i_2_5_98_0 & ~i_2_5_99_0) | (i_2_5_42_0 & ~i_2_5_90_0))) | (~i_2_5_65_0 & ((~i_2_5_90_0 & ~i_2_5_98_0) | (i_2_5_82_0 & (~i_2_5_99_0 | (i_2_5_42_0 & i_2_5_84_0 & ~i_2_5_90_0))))) | (i_2_5_42_0 & ((~i_2_5_98_0 & ~i_2_5_99_0) | (~i_2_5_90_0 & (~i_2_5_99_0 | (i_2_5_82_0 & ~i_2_5_98_0))))) | (~i_2_5_90_0 & ~i_2_5_98_0 & ~i_2_5_99_0))) | (i_2_5_42_0 & ((~i_2_5_65_0 & ((i_2_5_12_0 & ~i_2_5_98_0 & ~i_2_5_99_0) | (~i_2_5_90_0 & ((i_2_5_12_0 & (~i_2_5_99_0 | (i_2_5_82_0 & i_2_5_84_0))) | (~i_2_5_99_0 & (i_2_5_82_0 | i_2_5_84_0)))))) | (i_2_5_84_0 & ~i_2_5_90_0 & ~i_2_5_98_0 & ~i_2_5_99_0))) | (~i_2_5_65_0 & i_2_5_84_0 & ~i_2_5_98_0 & ~i_2_5_99_0))) | (~i_2_5_98_0 & ((~i_2_5_99_0 & ((i_2_5_12_0 & ((i_2_5_42_0 & (i_2_5_62_0 | (~i_2_5_65_0 & ~i_2_5_90_0))) | (~i_2_5_65_0 & i_2_5_82_0 & ~i_2_5_90_0) | (i_2_5_62_0 & ((i_2_5_82_0 & ~i_2_5_90_0) | ((~i_2_5_65_0 | i_2_5_84_0) & (i_2_5_82_0 | ~i_2_5_90_0)))))) | (~i_2_5_65_0 & ((i_2_5_42_0 & ((i_2_5_84_0 & ~i_2_5_90_0) | (~i_2_5_12_0 & i_2_5_82_0 & ~i_2_5_84_0))) | (i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_90_0) | (i_2_5_62_0 & ((i_2_5_84_0 & ~i_2_5_90_0) | (i_2_5_82_0 & (i_2_5_84_0 | ~i_2_5_90_0)))))) | (i_2_5_62_0 & i_2_5_84_0 & ~i_2_5_90_0 & (i_2_5_42_0 | i_2_5_82_0)))) | (~i_2_5_65_0 & i_2_5_84_0 & ((i_2_5_12_0 & (i_2_5_82_0 | (i_2_5_62_0 & i_2_5_90_0 & i_2_5_93_0))) | (i_2_5_42_0 & i_2_5_82_0 & ~i_2_5_90_0))))) | (~i_2_5_90_0 & ((i_2_5_62_0 & ((i_2_5_42_0 & ((~i_2_5_65_0 & i_2_5_84_0 & ~i_2_5_99_0) | (i_2_5_12_0 & (~i_2_5_99_0 | (i_2_5_84_0 & i_2_5_98_0))))) | (i_2_5_84_0 & ~i_2_5_99_0 & ~i_2_5_65_0 & i_2_5_82_0))) | (i_2_5_84_0 & ~i_2_5_99_0 & i_2_5_12_0 & ~i_2_5_65_0))))) | (i_2_5_62_0 & ((i_2_5_148_0 & ((~i_2_5_98_0 & ((i_2_5_12_0 & ((~i_2_5_90_0 & ~i_2_5_99_0) | (i_2_5_42_0 & ~i_2_5_84_0 & i_2_5_93_0 & ~i_2_5_102_0))) | (i_2_5_42_0 & ((~i_2_5_90_0 & ~i_2_5_99_0) | (~i_2_5_65_0 & i_2_5_84_0 & i_2_5_90_0 & i_2_5_93_0))) | (~i_2_5_99_0 & ((~i_2_5_65_0 & i_2_5_82_0 & i_2_5_84_0) | (i_2_5_65_0 & ~i_2_5_84_0 & ~i_2_5_90_0))))) | (~i_2_5_99_0 & ((i_2_5_82_0 & ~i_2_5_90_0 & (~i_2_5_65_0 | i_2_5_84_0)) | (i_2_5_12_0 & i_2_5_42_0 & i_2_5_90_0))))) | (~i_2_5_65_0 & ((i_2_5_84_0 & ((i_2_5_42_0 & ((i_2_5_82_0 & ~i_2_5_98_0) | (i_2_5_12_0 & ~i_2_5_148_0))) | (i_2_5_12_0 & ~i_2_5_99_0 & (i_2_5_82_0 | (~i_2_5_90_0 & ~i_2_5_98_0))) | (i_2_5_82_0 & ~i_2_5_90_0 & i_2_5_93_0 & ~i_2_5_98_0 & ~i_2_5_102_0 & ~i_2_5_148_0))) | (i_2_5_12_0 & i_2_5_82_0 & ~i_2_5_84_0 & ~i_2_5_90_0 & i_2_5_98_0 & ~i_2_5_148_0))))) | (i_2_5_12_0 & ((i_2_5_84_0 & ((~i_2_5_65_0 & ~i_2_5_98_0 & ((~i_2_5_99_0 & i_2_5_148_0) | (i_2_5_42_0 & (~i_2_5_90_0 | i_2_5_99_0)))) | (~i_2_5_99_0 & ((~i_2_5_90_0 & i_2_5_148_0) | (i_2_5_82_0 & (~i_2_5_90_0 | i_2_5_148_0)))))) | (i_2_5_42_0 & ~i_2_5_90_0 & ~i_2_5_98_0 & ~i_2_5_99_0 & i_2_5_148_0))) | (i_2_5_42_0 & ~i_2_5_65_0 & i_2_5_84_0 & ~i_2_5_99_0 & i_2_5_148_0 & ~i_2_5_90_0 & ~i_2_5_98_0))) | (~i_2_5_99_0 & ((~i_2_5_90_0 & ((i_2_5_62_0 & ((i_2_5_148_0 & ((i_2_5_42_0 & ((~i_2_5_65_0 & i_2_5_84_0) | (~i_2_5_82_0 & ~i_2_5_98_0 & i_2_5_102_0))) | (~i_2_5_42_0 & ((~i_2_5_65_0 & i_2_5_70_0 & ~i_2_5_98_0) | (i_2_5_82_0 & ~i_2_5_84_0 & i_2_5_93_0 & ~i_2_5_102_0))) | (i_2_5_102_0 & (i_2_5_12_0 | (i_2_5_84_0 & (~i_2_5_65_0 | (i_2_5_82_0 & ~i_2_5_98_0))))))) | (i_2_5_12_0 & ((~i_2_5_65_0 & ((i_2_5_82_0 & ~i_2_5_84_0) | (i_2_5_84_0 & ~i_2_5_98_0 & i_2_5_102_0))) | (i_2_5_42_0 & i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_98_0 & i_2_5_102_0))) | (~i_2_5_65_0 & i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_98_0 & i_2_5_102_0))) | (~i_2_5_65_0 & i_2_5_102_0 & ((~i_2_5_98_0 & ((i_2_5_42_0 & i_2_5_84_0 & i_2_5_148_0) | (i_2_5_12_0 & (i_2_5_148_0 | (i_2_5_82_0 & i_2_5_84_0))))) | (i_2_5_84_0 & i_2_5_148_0 & ~i_2_5_42_0 & i_2_5_82_0))) | (i_2_5_12_0 & i_2_5_82_0 & ~i_2_5_98_0 & ~i_2_5_102_0 & i_2_5_148_0))) | (i_2_5_62_0 & ((i_2_5_42_0 & i_2_5_102_0 & ((i_2_5_12_0 & ((i_2_5_84_0 & i_2_5_148_0) | (~i_2_5_65_0 & i_2_5_90_0 & ~i_2_5_98_0))) | (~i_2_5_65_0 & i_2_5_84_0 & ~i_2_5_98_0 & i_2_5_148_0))) | (i_2_5_82_0 & i_2_5_148_0 & i_2_5_12_0 & ~i_2_5_65_0))))) | (~i_2_5_65_0 & i_2_5_82_0 & ~i_2_5_98_0 & ((i_2_5_42_0 & i_2_5_62_0 & ((i_2_5_84_0 & i_2_5_102_0 & i_2_5_148_0) | (i_2_5_99_0 & ~i_2_5_148_0 & ~i_2_5_84_0 & ~i_2_5_90_0))) | (i_2_5_102_0 & i_2_5_148_0 & i_2_5_12_0 & ~i_2_5_90_0))))) | (i_2_5_102_0 & ((~i_2_5_98_0 & ((i_2_5_148_0 & ((~i_2_5_65_0 & ((~i_2_5_90_0 & ((~i_2_5_12_0 & ~i_2_5_84_0 & ((i_2_5_82_0 & i_2_5_93_0 & ~i_2_5_42_0 & i_2_5_62_0) | (~i_2_5_82_0 & ~i_2_5_99_0 & i_2_5_42_0 & ~i_2_5_70_0))) | (i_2_5_84_0 & ((i_2_5_62_0 & ((i_2_5_42_0 & ~i_2_5_99_0) | (~i_2_5_70_0 & i_2_5_82_0 & ~i_2_5_93_0))) | (~i_2_5_70_0 & i_2_5_82_0 & ~i_2_5_99_0) | (i_2_5_12_0 & i_2_5_70_0 & ~i_2_5_93_0))) | (i_2_5_82_0 & ~i_2_5_93_0 & ~i_2_5_99_0))) | (~i_2_5_99_0 & ((i_2_5_82_0 & ((i_2_5_62_0 & ((i_2_5_42_0 & ((i_2_5_12_0 & (i_2_5_84_0 | ~i_2_5_93_0)) | (i_2_5_84_0 & (~i_2_5_70_0 | ~i_2_5_93_0)))) | (~i_2_5_70_0 & ~i_2_5_93_0))) | (~i_2_5_70_0 & ~i_2_5_93_0 & (i_2_5_12_0 | i_2_5_84_0)))) | (i_2_5_12_0 & i_2_5_84_0 & (~i_2_5_70_0 | ~i_2_5_93_0)))) | (i_2_5_12_0 & i_2_5_62_0 & ~i_2_5_70_0 & i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_93_0))) | (~i_2_5_70_0 & ((i_2_5_62_0 & ((~i_2_5_99_0 & ((i_2_5_65_0 & ((i_2_5_12_0 & ~i_2_5_84_0 & i_2_5_93_0) | (~i_2_5_82_0 & ~i_2_5_93_0))) | (~i_2_5_93_0 & ((i_2_5_12_0 & ~i_2_5_82_0) | (i_2_5_42_0 & (~i_2_5_82_0 | i_2_5_84_0)))) | (i_2_5_12_0 & (~i_2_5_90_0 | (i_2_5_42_0 & i_2_5_82_0))))) | (i_2_5_42_0 & ~i_2_5_93_0 & ((~i_2_5_82_0 & i_2_5_84_0) | (i_2_5_82_0 & ~i_2_5_84_0 & ~i_2_5_90_0))))) | (i_2_5_12_0 & i_2_5_84_0 & ((~i_2_5_82_0 & ~i_2_5_99_0) | (~i_2_5_93_0 & (~i_2_5_99_0 | (i_2_5_65_0 & ~i_2_5_90_0))))))) | (i_2_5_12_0 & ~i_2_5_93_0 & ~i_2_5_99_0 & ((i_2_5_84_0 & (i_2_5_42_0 | ~i_2_5_90_0)) | (~i_2_5_42_0 & ~i_2_5_82_0 & ~i_2_5_90_0))))) | (~i_2_5_70_0 & ((~i_2_5_90_0 & ((i_2_5_42_0 & ((i_2_5_12_0 & ((i_2_5_82_0 & ~i_2_5_84_0 & i_2_5_92_0 & ~i_2_5_93_0) | (i_2_5_62_0 & i_2_5_84_0 & ~i_2_5_99_0))) | (i_2_5_62_0 & ~i_2_5_99_0 & ((i_2_5_84_0 & ~i_2_5_93_0) | (~i_2_5_65_0 & (i_2_5_82_0 | ~i_2_5_84_0)))))) | (~i_2_5_65_0 & ((i_2_5_82_0 & ((i_2_5_12_0 & i_2_5_84_0 & (~i_2_5_99_0 | (i_2_5_62_0 & ~i_2_5_93_0))) | (i_2_5_62_0 & ~i_2_5_93_0 & ~i_2_5_99_0))) | (i_2_5_62_0 & i_2_5_84_0 & ~i_2_5_93_0 & ~i_2_5_99_0))) | (i_2_5_12_0 & i_2_5_84_0 & ~i_2_5_93_0 & ~i_2_5_99_0))) | (i_2_5_62_0 & ~i_2_5_65_0 & ~i_2_5_99_0 & ((i_2_5_12_0 & ((i_2_5_84_0 & ~i_2_5_93_0) | (i_2_5_42_0 & i_2_5_82_0 & (i_2_5_84_0 | ~i_2_5_93_0)))) | (i_2_5_42_0 & i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_93_0))))))) | (~i_2_5_99_0 & ((~i_2_5_93_0 & ((i_2_5_62_0 & ((~i_2_5_65_0 & ((i_2_5_42_0 & ((i_2_5_12_0 & i_2_5_84_0) | (i_2_5_70_0 & i_2_5_82_0 & ~i_2_5_90_0))) | (~i_2_5_70_0 & ((i_2_5_12_0 & (~i_2_5_90_0 | (i_2_5_82_0 & i_2_5_148_0))) | (i_2_5_148_0 & (~i_2_5_90_0 | (i_2_5_82_0 & i_2_5_84_0))))) | (i_2_5_84_0 & ((i_2_5_12_0 & ~i_2_5_90_0) | (~i_2_5_42_0 & ~i_2_5_82_0 & i_2_5_148_0))))) | (~i_2_5_90_0 & i_2_5_148_0 & ~i_2_5_42_0 & ~i_2_5_70_0))) | (i_2_5_84_0 & ((i_2_5_12_0 & i_2_5_42_0 & (~i_2_5_70_0 | (i_2_5_82_0 & ~i_2_5_90_0))) | (~i_2_5_70_0 & i_2_5_82_0 & ~i_2_5_90_0 & (~i_2_5_65_0 | i_2_5_148_0)))) | (~i_2_5_90_0 & i_2_5_148_0 & i_2_5_12_0 & ~i_2_5_70_0))) | (i_2_5_42_0 & i_2_5_62_0 & ((~i_2_5_65_0 & ((i_2_5_12_0 & i_2_5_82_0 & (~i_2_5_90_0 | (~i_2_5_70_0 & i_2_5_84_0 & i_2_5_148_0))) | (~i_2_5_90_0 & i_2_5_148_0 & ~i_2_5_70_0 & i_2_5_84_0))) | (~i_2_5_70_0 & ~i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_90_0 & i_2_5_148_0))) | (i_2_5_82_0 & ~i_2_5_90_0 & i_2_5_148_0 & i_2_5_12_0 & ~i_2_5_70_0))) | (i_2_5_62_0 & ~i_2_5_65_0 & ~i_2_5_70_0 & ~i_2_5_90_0 & ((i_2_5_12_0 & i_2_5_84_0 & (i_2_5_42_0 | i_2_5_148_0)) | (i_2_5_42_0 & i_2_5_82_0 & ~i_2_5_84_0 & i_2_5_93_0 & i_2_5_99_0 & ~i_2_5_148_0))))) | (i_2_5_62_0 & ((~i_2_5_93_0 & ((~i_2_5_99_0 & ((i_2_5_148_0 & ((~i_2_5_70_0 & ((i_2_5_82_0 & ((~i_2_5_42_0 & ~i_2_5_90_0) | (~i_2_5_65_0 & ((i_2_5_84_0 & ~i_2_5_98_0) | (i_2_5_12_0 & (~i_2_5_42_0 | ~i_2_5_98_0)))))) | (~i_2_5_65_0 & ~i_2_5_98_0 & ((i_2_5_12_0 & i_2_5_84_0) | (i_2_5_42_0 & ~i_2_5_90_0))))) | (i_2_5_12_0 & ((~i_2_5_65_0 & (~i_2_5_90_0 | (i_2_5_42_0 & i_2_5_82_0 & i_2_5_84_0))) | (i_2_5_42_0 & (~i_2_5_90_0 | (i_2_5_84_0 & ~i_2_5_102_0 & i_2_5_65_0 & i_2_5_70_0))))) | (i_2_5_42_0 & i_2_5_82_0 & i_2_5_84_0 & ~i_2_5_90_0 & ~i_2_5_98_0))) | (~i_2_5_65_0 & ~i_2_5_70_0 & ~i_2_5_90_0 & ~i_2_5_98_0 & ((i_2_5_42_0 & i_2_5_82_0) | (i_2_5_12_0 & i_2_5_84_0))))) | (i_2_5_12_0 & i_2_5_42_0 & ~i_2_5_65_0 & ~i_2_5_70_0 & ~i_2_5_98_0 & (~i_2_5_90_0 | (~i_2_5_102_0 & ~i_2_5_148_0 & i_2_5_82_0 & i_2_5_84_0))))) | (~i_2_5_70_0 & ~i_2_5_98_0 & ~i_2_5_99_0 & ((i_2_5_12_0 & i_2_5_42_0 & ((~i_2_5_65_0 & ~i_2_5_90_0 & ~i_2_5_148_0) | (i_2_5_82_0 & i_2_5_84_0 & i_2_5_148_0))) | (i_2_5_84_0 & ~i_2_5_90_0 & i_2_5_148_0 & ~i_2_5_42_0 & ~i_2_5_65_0))))) | (i_2_5_12_0 & ~i_2_5_93_0 & ((~i_2_5_98_0 & i_2_5_148_0 & ((i_2_5_82_0 & ~i_2_5_90_0 & ~i_2_5_42_0 & ~i_2_5_65_0) | (i_2_5_84_0 & ~i_2_5_99_0 & i_2_5_42_0 & ~i_2_5_70_0))) | (i_2_5_82_0 & ~i_2_5_90_0 & ~i_2_5_99_0 & ((~i_2_5_65_0 & ~i_2_5_70_0) | (i_2_5_42_0 & ~i_2_5_102_0 & (~i_2_5_65_0 | ~i_2_5_70_0))))));
endmodule
