module ee681proj4 ( 
    i_2_0_13_0, i_2_0_16_0, i_2_0_49_0, i_2_0_57_0, i_2_0_66_0, i_2_0_74_0,
    i_2_0_78_0, i_2_0_94_0, i_2_0_97_0, i_2_0_109_0, i_2_0_118_0,
    i_2_0_139_0, i_2_0_142_0, i_2_0_143_0, i_2_0_147_0,
    o_2_0_0_0  );
  input  i_2_0_13_0, i_2_0_16_0, i_2_0_49_0, i_2_0_57_0, i_2_0_66_0,
    i_2_0_74_0, i_2_0_78_0, i_2_0_94_0, i_2_0_97_0, i_2_0_109_0,
    i_2_0_118_0, i_2_0_139_0, i_2_0_142_0, i_2_0_143_0, i_2_0_147_0;
  output o_2_0_0_0;
  wire new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_;
  NOT      g0000(.a(i_2_0_143_0), .O(new_n17_));
  NOT      g0001(.a(i_2_0_94_0), .O(new_n18_));
  OR       g0002(.a(i_2_0_109_0), .b(i_2_0_78_0), .O(new_n19_));
  NOT      g0003(.a(new_n19_), .O(new_n20_));
  NOT      g0004(.a(i_2_0_139_0), .O(new_n21_));
  AND      g0005(.a(new_n21_), .b(i_2_0_16_0), .O(new_n22_));
  NOT      g0006(.a(i_2_0_97_0), .O(new_n23_));
  NOT      g0007(.a(i_2_0_147_0), .O(new_n24_));
  AND      g0008(.a(new_n24_), .b(i_2_0_118_0), .O(new_n25_));
  OR       g0009(.a(new_n25_), .b(new_n23_), .O(new_n26_));
  AND      g0010(.a(new_n26_), .b(new_n22_), .O(new_n27_));
  OR       g0011(.a(i_2_0_147_0), .b(i_2_0_142_0), .O(new_n28_));
  NOT      g0012(.a(i_2_0_118_0), .O(new_n29_));
  AND      g0013(.a(i_2_0_97_0), .b(i_2_0_74_0), .O(new_n30_));
  AND      g0014(.a(new_n30_), .b(new_n29_), .O(new_n31_));
  OR       g0015(.a(new_n31_), .b(new_n28_), .O(new_n32_));
  NOT      g0016(.a(i_2_0_74_0), .O(new_n33_));
  AND      g0017(.a(new_n33_), .b(i_2_0_16_0), .O(new_n34_));
  OR       g0018(.a(i_2_0_147_0), .b(i_2_0_97_0), .O(new_n35_));
  NAND     g0019(.a(new_n35_), .b(new_n29_), .O(new_n36_));
  NAND     g0020(.a(new_n36_), .b(new_n34_), .O(new_n37_));
  NAND     g0021(.a(new_n37_), .b(new_n32_), .O(new_n38_));
  OR       g0022(.a(new_n38_), .b(new_n27_), .O(new_n39_));
  AND      g0023(.a(new_n39_), .b(new_n20_), .O(new_n40_));
  NOT      g0024(.a(i_2_0_16_0), .O(new_n41_));
  OR       g0025(.a(i_2_0_139_0), .b(new_n29_), .O(new_n42_));
  OR       g0026(.a(new_n42_), .b(new_n41_), .O(new_n43_));
  OR       g0027(.a(i_2_0_142_0), .b(new_n41_), .O(new_n44_));
  OR       g0028(.a(i_2_0_142_0), .b(i_2_0_139_0), .O(new_n45_));
  AND      g0029(.a(new_n45_), .b(new_n44_), .O(new_n46_));
  NAND     g0030(.a(new_n46_), .b(new_n43_), .O(new_n47_));
  AND      g0031(.a(i_2_0_147_0), .b(i_2_0_109_0), .O(new_n48_));
  OR       g0032(.a(new_n48_), .b(i_2_0_142_0), .O(new_n49_));
  NAND     g0033(.a(new_n49_), .b(i_2_0_74_0), .O(new_n50_));
  OR       g0034(.a(i_2_0_147_0), .b(i_2_0_109_0), .O(new_n51_));
  AND      g0035(.a(new_n51_), .b(i_2_0_142_0), .O(new_n52_));
  OR       g0036(.a(new_n52_), .b(i_2_0_57_0), .O(new_n53_));
  OR       g0037(.a(i_2_0_142_0), .b(i_2_0_74_0), .O(new_n54_));
  OR       g0038(.a(new_n54_), .b(new_n48_), .O(new_n55_));
  NAND     g0039(.a(new_n55_), .b(new_n53_), .O(new_n56_));
  AND      g0040(.a(new_n56_), .b(new_n50_), .O(new_n57_));
  OR       g0041(.a(new_n57_), .b(new_n47_), .O(new_n58_));
  AND      g0042(.a(new_n58_), .b(new_n23_), .O(new_n59_));
  OR       g0043(.a(new_n59_), .b(new_n40_), .O(new_n60_));
  NAND     g0044(.a(i_2_0_139_0), .b(i_2_0_109_0), .O(new_n61_));
  NOT      g0045(.a(i_2_0_78_0), .O(new_n62_));
  NOT      g0046(.a(i_2_0_57_0), .O(new_n63_));
  AND      g0047(.a(new_n63_), .b(i_2_0_16_0), .O(new_n64_));
  AND      g0048(.a(new_n64_), .b(new_n62_), .O(new_n65_));
  AND      g0049(.a(new_n65_), .b(new_n61_), .O(new_n66_));
  OR       g0050(.a(i_2_0_142_0), .b(i_2_0_78_0), .O(new_n67_));
  NOT      g0051(.a(new_n67_), .O(new_n68_));
  NAND     g0052(.a(i_2_0_139_0), .b(i_2_0_74_0), .O(new_n69_));
  NAND     g0053(.a(new_n69_), .b(i_2_0_118_0), .O(new_n70_));
  OR       g0054(.a(new_n48_), .b(i_2_0_139_0), .O(new_n71_));
  NAND     g0055(.a(new_n71_), .b(new_n70_), .O(new_n72_));
  AND      g0056(.a(new_n72_), .b(new_n68_), .O(new_n73_));
  OR       g0057(.a(new_n73_), .b(new_n66_), .O(new_n74_));
  OR       g0058(.a(i_2_0_78_0), .b(i_2_0_57_0), .O(new_n75_));
  NOT      g0059(.a(new_n75_), .O(new_n76_));
  OR       g0060(.a(i_2_0_139_0), .b(i_2_0_74_0), .O(new_n77_));
  OR       g0061(.a(new_n29_), .b(i_2_0_109_0), .O(new_n78_));
  OR       g0062(.a(new_n78_), .b(i_2_0_147_0), .O(new_n79_));
  AND      g0063(.a(new_n79_), .b(new_n35_), .O(new_n80_));
  OR       g0064(.a(new_n80_), .b(new_n77_), .O(new_n81_));
  NOT      g0065(.a(i_2_0_142_0), .O(new_n82_));
  NOT      g0066(.a(new_n48_), .O(new_n83_));
  OR       g0067(.a(i_2_0_118_0), .b(new_n33_), .O(new_n84_));
  OR       g0068(.a(new_n84_), .b(new_n83_), .O(new_n85_));
  NAND     g0069(.a(new_n85_), .b(new_n82_), .O(new_n86_));
  NAND     g0070(.a(new_n86_), .b(new_n81_), .O(new_n87_));
  AND      g0071(.a(new_n87_), .b(new_n76_), .O(new_n88_));
  OR       g0072(.a(new_n88_), .b(new_n74_), .O(new_n89_));
  OR       g0073(.a(new_n89_), .b(new_n60_), .O(new_n90_));
  OR       g0074(.a(new_n24_), .b(i_2_0_118_0), .O(new_n91_));
  OR       g0075(.a(i_2_0_74_0), .b(i_2_0_57_0), .O(new_n92_));
  NAND     g0076(.a(new_n92_), .b(new_n41_), .O(new_n93_));
  AND      g0077(.a(new_n93_), .b(new_n91_), .O(new_n94_));
  AND      g0078(.a(i_2_0_74_0), .b(i_2_0_57_0), .O(new_n95_));
  OR       g0079(.a(new_n95_), .b(i_2_0_139_0), .O(new_n96_));
  OR       g0080(.a(i_2_0_147_0), .b(new_n29_), .O(new_n97_));
  AND      g0081(.a(i_2_0_139_0), .b(i_2_0_57_0), .O(new_n98_));
  OR       g0082(.a(new_n98_), .b(new_n97_), .O(new_n99_));
  NAND     g0083(.a(new_n99_), .b(new_n96_), .O(new_n100_));
  OR       g0084(.a(new_n100_), .b(new_n94_), .O(new_n101_));
  AND      g0085(.a(new_n101_), .b(new_n82_), .O(new_n102_));
  OR       g0086(.a(new_n95_), .b(i_2_0_109_0), .O(new_n103_));
  OR       g0087(.a(i_2_0_139_0), .b(new_n41_), .O(new_n104_));
  OR       g0088(.a(i_2_0_142_0), .b(new_n29_), .O(new_n105_));
  NAND     g0089(.a(new_n105_), .b(new_n104_), .O(new_n106_));
  NAND     g0090(.a(i_2_0_147_0), .b(i_2_0_57_0), .O(new_n107_));
  NAND     g0091(.a(new_n107_), .b(new_n106_), .O(new_n108_));
  OR       g0092(.a(new_n108_), .b(new_n103_), .O(new_n109_));
  OR       g0093(.a(i_2_0_142_0), .b(i_2_0_109_0), .O(new_n110_));
  NOT      g0094(.a(new_n110_), .O(new_n111_));
  AND      g0095(.a(new_n91_), .b(new_n21_), .O(new_n112_));
  OR       g0096(.a(i_2_0_147_0), .b(i_2_0_57_0), .O(new_n113_));
  NOT      g0097(.a(new_n113_), .O(new_n114_));
  OR       g0098(.a(new_n114_), .b(new_n93_), .O(new_n115_));
  OR       g0099(.a(new_n115_), .b(new_n112_), .O(new_n116_));
  NAND     g0100(.a(new_n116_), .b(new_n111_), .O(new_n117_));
  NAND     g0101(.a(new_n117_), .b(new_n109_), .O(new_n118_));
  OR       g0102(.a(new_n118_), .b(new_n102_), .O(new_n119_));
  OR       g0103(.a(new_n42_), .b(new_n62_), .O(new_n120_));
  OR       g0104(.a(i_2_0_74_0), .b(new_n63_), .O(new_n121_));
  OR       g0105(.a(new_n121_), .b(new_n120_), .O(new_n122_));
  OR       g0106(.a(new_n21_), .b(i_2_0_118_0), .O(new_n123_));
  OR       g0107(.a(i_2_0_97_0), .b(i_2_0_78_0), .O(new_n124_));
  OR       g0108(.a(new_n124_), .b(new_n92_), .O(new_n125_));
  NAND     g0109(.a(i_2_0_78_0), .b(i_2_0_16_0), .O(new_n126_));
  OR       g0110(.a(new_n126_), .b(i_2_0_57_0), .O(new_n127_));
  AND      g0111(.a(new_n127_), .b(new_n125_), .O(new_n128_));
  OR       g0112(.a(new_n128_), .b(new_n123_), .O(new_n129_));
  NAND     g0113(.a(new_n129_), .b(new_n122_), .O(new_n130_));
  AND      g0114(.a(new_n130_), .b(i_2_0_147_0), .O(new_n131_));
  NOT      g0115(.a(new_n124_), .O(new_n132_));
  AND      g0116(.a(new_n106_), .b(new_n24_), .O(new_n133_));
  AND      g0117(.a(new_n24_), .b(i_2_0_16_0), .O(new_n134_));
  AND      g0118(.a(i_2_0_118_0), .b(i_2_0_109_0), .O(new_n135_));
  AND      g0119(.a(new_n135_), .b(new_n134_), .O(new_n136_));
  OR       g0120(.a(i_2_0_139_0), .b(i_2_0_109_0), .O(new_n137_));
  OR       g0121(.a(new_n29_), .b(i_2_0_57_0), .O(new_n138_));
  OR       g0122(.a(new_n138_), .b(new_n137_), .O(new_n139_));
  OR       g0123(.a(new_n95_), .b(i_2_0_142_0), .O(new_n140_));
  NAND     g0124(.a(new_n140_), .b(new_n139_), .O(new_n141_));
  OR       g0125(.a(new_n141_), .b(new_n136_), .O(new_n142_));
  OR       g0126(.a(new_n142_), .b(new_n133_), .O(new_n143_));
  AND      g0127(.a(new_n143_), .b(new_n132_), .O(new_n144_));
  OR       g0128(.a(new_n144_), .b(new_n131_), .O(new_n145_));
  OR       g0129(.a(new_n145_), .b(new_n119_), .O(new_n146_));
  OR       g0130(.a(new_n146_), .b(new_n90_), .O(new_n147_));
  AND      g0131(.a(new_n147_), .b(i_2_0_13_0), .O(new_n148_));
  AND      g0132(.a(new_n82_), .b(i_2_0_16_0), .O(new_n149_));
  OR       g0133(.a(i_2_0_139_0), .b(i_2_0_78_0), .O(new_n150_));
  NOT      g0134(.a(new_n150_), .O(new_n151_));
  NOT      g0135(.a(i_2_0_109_0), .O(new_n152_));
  OR       g0136(.a(i_2_0_118_0), .b(new_n152_), .O(new_n153_));
  NAND     g0137(.a(i_2_0_139_0), .b(i_2_0_78_0), .O(new_n154_));
  AND      g0138(.a(new_n154_), .b(new_n153_), .O(new_n155_));
  OR       g0139(.a(i_2_0_147_0), .b(i_2_0_139_0), .O(new_n156_));
  NAND     g0140(.a(new_n79_), .b(new_n156_), .O(new_n157_));
  OR       g0141(.a(new_n157_), .b(new_n155_), .O(new_n158_));
  OR       g0142(.a(new_n24_), .b(i_2_0_78_0), .O(new_n159_));
  AND      g0143(.a(new_n159_), .b(new_n158_), .O(new_n160_));
  OR       g0144(.a(new_n160_), .b(new_n151_), .O(new_n161_));
  AND      g0145(.a(new_n161_), .b(new_n23_), .O(new_n162_));
  NOT      g0146(.a(new_n98_), .O(new_n163_));
  OR       g0147(.a(i_2_0_118_0), .b(new_n62_), .O(new_n164_));
  NAND     g0148(.a(new_n156_), .b(i_2_0_109_0), .O(new_n165_));
  AND      g0149(.a(new_n165_), .b(new_n164_), .O(new_n166_));
  AND      g0150(.a(new_n166_), .b(new_n163_), .O(new_n167_));
  OR       g0151(.a(i_2_0_78_0), .b(i_2_0_74_0), .O(new_n168_));
  NOT      g0152(.a(new_n168_), .O(new_n169_));
  AND      g0153(.a(i_2_0_118_0), .b(new_n62_), .O(new_n170_));
  OR       g0154(.a(new_n170_), .b(new_n169_), .O(new_n171_));
  AND      g0155(.a(new_n51_), .b(i_2_0_57_0), .O(new_n172_));
  NAND     g0156(.a(new_n172_), .b(new_n70_), .O(new_n173_));
  AND      g0157(.a(new_n173_), .b(new_n171_), .O(new_n174_));
  OR       g0158(.a(i_2_0_147_0), .b(new_n152_), .O(new_n175_));
  AND      g0159(.a(i_2_0_118_0), .b(new_n33_), .O(new_n176_));
  NOT      g0160(.a(new_n156_), .O(new_n177_));
  OR       g0161(.a(new_n177_), .b(new_n176_), .O(new_n178_));
  AND      g0162(.a(new_n178_), .b(new_n175_), .O(new_n179_));
  OR       g0163(.a(new_n113_), .b(i_2_0_78_0), .O(new_n180_));
  NAND     g0164(.a(new_n180_), .b(new_n96_), .O(new_n181_));
  OR       g0165(.a(new_n181_), .b(new_n179_), .O(new_n182_));
  OR       g0166(.a(new_n182_), .b(new_n174_), .O(new_n183_));
  OR       g0167(.a(new_n183_), .b(new_n167_), .O(new_n184_));
  OR       g0168(.a(new_n184_), .b(new_n162_), .O(new_n185_));
  AND      g0169(.a(new_n185_), .b(new_n149_), .O(new_n186_));
  AND      g0170(.a(new_n23_), .b(i_2_0_16_0), .O(new_n187_));
  OR       g0171(.a(i_2_0_142_0), .b(i_2_0_57_0), .O(new_n188_));
  OR       g0172(.a(i_2_0_147_0), .b(i_2_0_78_0), .O(new_n189_));
  OR       g0173(.a(new_n189_), .b(new_n139_), .O(new_n190_));
  AND      g0174(.a(new_n190_), .b(new_n188_), .O(new_n191_));
  AND      g0175(.a(new_n48_), .b(i_2_0_57_0), .O(new_n192_));
  NAND     g0176(.a(new_n150_), .b(new_n29_), .O(new_n193_));
  AND      g0177(.a(new_n193_), .b(new_n192_), .O(new_n194_));
  AND      g0178(.a(new_n29_), .b(i_2_0_57_0), .O(new_n195_));
  OR       g0179(.a(new_n19_), .b(i_2_0_139_0), .O(new_n196_));
  OR       g0180(.a(new_n196_), .b(new_n195_), .O(new_n197_));
  AND      g0181(.a(new_n49_), .b(new_n67_), .O(new_n198_));
  NAND     g0182(.a(new_n198_), .b(new_n197_), .O(new_n199_));
  OR       g0183(.a(new_n199_), .b(new_n194_), .O(new_n200_));
  NAND     g0184(.a(new_n200_), .b(new_n33_), .O(new_n201_));
  NAND     g0185(.a(new_n201_), .b(new_n191_), .O(new_n202_));
  AND      g0186(.a(new_n202_), .b(new_n187_), .O(new_n203_));
  NOT      g0187(.a(new_n45_), .O(new_n204_));
  OR       g0188(.a(new_n97_), .b(new_n92_), .O(new_n205_));
  OR       g0189(.a(new_n78_), .b(new_n113_), .O(new_n206_));
  OR       g0190(.a(i_2_0_97_0), .b(i_2_0_74_0), .O(new_n207_));
  OR       g0191(.a(new_n207_), .b(new_n51_), .O(new_n208_));
  AND      g0192(.a(new_n208_), .b(new_n206_), .O(new_n209_));
  NAND     g0193(.a(new_n209_), .b(new_n205_), .O(new_n210_));
  OR       g0194(.a(new_n29_), .b(i_2_0_78_0), .O(new_n211_));
  AND      g0195(.a(new_n211_), .b(i_2_0_57_0), .O(new_n212_));
  AND      g0196(.a(new_n207_), .b(new_n51_), .O(new_n213_));
  OR       g0197(.a(new_n213_), .b(new_n30_), .O(new_n214_));
  OR       g0198(.a(new_n214_), .b(new_n212_), .O(new_n215_));
  AND      g0199(.a(new_n207_), .b(new_n75_), .O(new_n216_));
  OR       g0200(.a(new_n216_), .b(new_n48_), .O(new_n217_));
  OR       g0201(.a(new_n30_), .b(i_2_0_78_0), .O(new_n218_));
  AND      g0202(.a(new_n218_), .b(new_n29_), .O(new_n219_));
  OR       g0203(.a(new_n219_), .b(new_n217_), .O(new_n220_));
  NAND     g0204(.a(new_n220_), .b(new_n215_), .O(new_n221_));
  OR       g0205(.a(new_n221_), .b(new_n210_), .O(new_n222_));
  AND      g0206(.a(new_n222_), .b(new_n204_), .O(new_n223_));
  NAND     g0207(.a(i_2_0_147_0), .b(i_2_0_118_0), .O(new_n224_));
  OR       g0208(.a(new_n224_), .b(i_2_0_57_0), .O(new_n225_));
  OR       g0209(.a(new_n48_), .b(i_2_0_74_0), .O(new_n226_));
  NAND     g0210(.a(new_n226_), .b(new_n225_), .O(new_n227_));
  OR       g0211(.a(i_2_0_142_0), .b(i_2_0_97_0), .O(new_n228_));
  NOT      g0212(.a(new_n228_), .O(new_n229_));
  AND      g0213(.a(i_2_0_118_0), .b(new_n152_), .O(new_n230_));
  OR       g0214(.a(new_n230_), .b(new_n63_), .O(new_n231_));
  AND      g0215(.a(new_n231_), .b(new_n62_), .O(new_n232_));
  AND      g0216(.a(new_n232_), .b(new_n229_), .O(new_n233_));
  AND      g0217(.a(new_n233_), .b(new_n227_), .O(new_n234_));
  OR       g0218(.a(new_n234_), .b(new_n223_), .O(new_n235_));
  OR       g0219(.a(new_n235_), .b(new_n203_), .O(new_n236_));
  OR       g0220(.a(new_n236_), .b(new_n186_), .O(new_n237_));
  OR       g0221(.a(new_n237_), .b(new_n148_), .O(new_n238_));
  AND      g0222(.a(new_n238_), .b(i_2_0_66_0), .O(new_n239_));
  AND      g0223(.a(new_n123_), .b(new_n23_), .O(new_n240_));
  NAND     g0224(.a(new_n240_), .b(new_n61_), .O(new_n241_));
  NAND     g0225(.a(new_n241_), .b(new_n120_), .O(new_n242_));
  AND      g0226(.a(new_n242_), .b(i_2_0_13_0), .O(new_n243_));
  OR       g0227(.a(new_n243_), .b(new_n82_), .O(new_n244_));
  AND      g0228(.a(i_2_0_139_0), .b(new_n62_), .O(new_n245_));
  OR       g0229(.a(new_n245_), .b(new_n97_), .O(new_n246_));
  NOT      g0230(.a(i_2_0_13_0), .O(new_n247_));
  OR       g0231(.a(i_2_0_109_0), .b(new_n23_), .O(new_n248_));
  AND      g0232(.a(new_n248_), .b(new_n247_), .O(new_n249_));
  OR       g0233(.a(new_n249_), .b(i_2_0_147_0), .O(new_n250_));
  NAND     g0234(.a(new_n250_), .b(new_n246_), .O(new_n251_));
  AND      g0235(.a(new_n251_), .b(new_n244_), .O(new_n252_));
  NAND     g0236(.a(i_2_0_142_0), .b(i_2_0_109_0), .O(new_n253_));
  OR       g0237(.a(new_n253_), .b(new_n166_), .O(new_n254_));
  OR       g0238(.a(new_n124_), .b(new_n29_), .O(new_n255_));
  OR       g0239(.a(new_n156_), .b(i_2_0_97_0), .O(new_n256_));
  AND      g0240(.a(new_n256_), .b(new_n228_), .O(new_n257_));
  NAND     g0241(.a(new_n257_), .b(new_n255_), .O(new_n258_));
  AND      g0242(.a(new_n258_), .b(new_n254_), .O(new_n259_));
  AND      g0243(.a(new_n21_), .b(i_2_0_97_0), .O(new_n260_));
  AND      g0244(.a(new_n29_), .b(i_2_0_109_0), .O(new_n261_));
  AND      g0245(.a(new_n261_), .b(i_2_0_13_0), .O(new_n262_));
  AND      g0246(.a(new_n262_), .b(new_n260_), .O(new_n263_));
  NOT      g0247(.a(new_n28_), .O(new_n264_));
  AND      g0248(.a(new_n264_), .b(i_2_0_78_0), .O(new_n265_));
  OR       g0249(.a(new_n265_), .b(new_n263_), .O(new_n266_));
  OR       g0250(.a(new_n266_), .b(new_n259_), .O(new_n267_));
  AND      g0251(.a(new_n267_), .b(new_n33_), .O(new_n268_));
  NAND     g0252(.a(new_n42_), .b(new_n247_), .O(new_n269_));
  AND      g0253(.a(new_n269_), .b(new_n111_), .O(new_n270_));
  OR       g0254(.a(new_n270_), .b(new_n268_), .O(new_n271_));
  OR       g0255(.a(new_n271_), .b(new_n252_), .O(new_n272_));
  AND      g0256(.a(new_n272_), .b(new_n64_), .O(new_n273_));
  AND      g0257(.a(new_n207_), .b(new_n70_), .O(new_n274_));
  NAND     g0258(.a(new_n274_), .b(new_n218_), .O(new_n275_));
  AND      g0259(.a(new_n275_), .b(i_2_0_13_0), .O(new_n276_));
  OR       g0260(.a(new_n42_), .b(i_2_0_78_0), .O(new_n277_));
  NAND     g0261(.a(new_n277_), .b(new_n77_), .O(new_n278_));
  AND      g0262(.a(new_n164_), .b(new_n23_), .O(new_n279_));
  AND      g0263(.a(new_n279_), .b(new_n278_), .O(new_n280_));
  OR       g0264(.a(new_n280_), .b(new_n276_), .O(new_n281_));
  AND      g0265(.a(new_n281_), .b(new_n83_), .O(new_n282_));
  NOT      g0266(.a(new_n51_), .O(new_n283_));
  NOT      g0267(.a(new_n30_), .O(new_n284_));
  OR       g0268(.a(new_n269_), .b(new_n151_), .O(new_n285_));
  AND      g0269(.a(new_n285_), .b(new_n284_), .O(new_n286_));
  OR       g0270(.a(new_n77_), .b(i_2_0_97_0), .O(new_n287_));
  NAND     g0271(.a(new_n287_), .b(new_n247_), .O(new_n288_));
  OR       g0272(.a(new_n170_), .b(new_n21_), .O(new_n289_));
  AND      g0273(.a(new_n289_), .b(new_n288_), .O(new_n290_));
  OR       g0274(.a(new_n290_), .b(new_n286_), .O(new_n291_));
  AND      g0275(.a(new_n291_), .b(new_n283_), .O(new_n292_));
  OR       g0276(.a(i_2_0_97_0), .b(new_n247_), .O(new_n293_));
  NOT      g0277(.a(new_n293_), .O(new_n294_));
  AND      g0278(.a(new_n294_), .b(new_n123_), .O(new_n295_));
  NOT      g0279(.a(new_n196_), .O(new_n296_));
  OR       g0280(.a(new_n176_), .b(i_2_0_13_0), .O(new_n297_));
  AND      g0281(.a(new_n297_), .b(new_n296_), .O(new_n298_));
  OR       g0282(.a(new_n298_), .b(new_n295_), .O(new_n299_));
  OR       g0283(.a(new_n299_), .b(new_n292_), .O(new_n300_));
  OR       g0284(.a(new_n300_), .b(new_n282_), .O(new_n301_));
  AND      g0285(.a(new_n301_), .b(new_n149_), .O(new_n302_));
  NOT      g0286(.a(new_n188_), .O(new_n303_));
  NOT      g0287(.a(new_n207_), .O(new_n304_));
  AND      g0288(.a(new_n152_), .b(i_2_0_13_0), .O(new_n305_));
  OR       g0289(.a(new_n305_), .b(new_n24_), .O(new_n306_));
  OR       g0290(.a(i_2_0_118_0), .b(i_2_0_13_0), .O(new_n307_));
  NAND     g0291(.a(new_n307_), .b(new_n62_), .O(new_n308_));
  NAND     g0292(.a(new_n308_), .b(new_n196_), .O(new_n309_));
  AND      g0293(.a(new_n309_), .b(new_n306_), .O(new_n310_));
  AND      g0294(.a(new_n24_), .b(i_2_0_139_0), .O(new_n311_));
  OR       g0295(.a(new_n311_), .b(new_n261_), .O(new_n312_));
  OR       g0296(.a(new_n61_), .b(i_2_0_118_0), .O(new_n313_));
  OR       g0297(.a(i_2_0_118_0), .b(i_2_0_78_0), .O(new_n314_));
  AND      g0298(.a(new_n314_), .b(new_n313_), .O(new_n315_));
  AND      g0299(.a(new_n315_), .b(new_n312_), .O(new_n316_));
  OR       g0300(.a(new_n316_), .b(new_n310_), .O(new_n317_));
  AND      g0301(.a(new_n317_), .b(new_n304_), .O(new_n318_));
  OR       g0302(.a(new_n78_), .b(new_n21_), .O(new_n319_));
  OR       g0303(.a(new_n319_), .b(new_n124_), .O(new_n320_));
  NOT      g0304(.a(new_n77_), .O(new_n321_));
  AND      g0305(.a(new_n321_), .b(i_2_0_13_0), .O(new_n322_));
  AND      g0306(.a(new_n169_), .b(new_n25_), .O(new_n323_));
  AND      g0307(.a(new_n323_), .b(i_2_0_139_0), .O(new_n324_));
  OR       g0308(.a(new_n324_), .b(new_n322_), .O(new_n325_));
  AND      g0309(.a(new_n193_), .b(i_2_0_13_0), .O(new_n326_));
  OR       g0310(.a(new_n326_), .b(new_n152_), .O(new_n327_));
  NAND     g0311(.a(new_n327_), .b(new_n325_), .O(new_n328_));
  NAND     g0312(.a(new_n328_), .b(new_n320_), .O(new_n329_));
  OR       g0313(.a(new_n329_), .b(new_n318_), .O(new_n330_));
  AND      g0314(.a(new_n330_), .b(new_n303_), .O(new_n331_));
  AND      g0315(.a(new_n279_), .b(new_n283_), .O(new_n332_));
  NOT      g0316(.a(new_n189_), .O(new_n333_));
  AND      g0317(.a(new_n333_), .b(new_n153_), .O(new_n334_));
  OR       g0318(.a(new_n230_), .b(new_n23_), .O(new_n335_));
  NAND     g0319(.a(i_2_0_147_0), .b(i_2_0_78_0), .O(new_n336_));
  AND      g0320(.a(new_n336_), .b(new_n335_), .O(new_n337_));
  OR       g0321(.a(new_n337_), .b(new_n334_), .O(new_n338_));
  NOT      g0322(.a(new_n95_), .O(new_n339_));
  NAND     g0323(.a(new_n189_), .b(i_2_0_109_0), .O(new_n340_));
  OR       g0324(.a(new_n340_), .b(new_n63_), .O(new_n341_));
  AND      g0325(.a(new_n341_), .b(new_n339_), .O(new_n342_));
  AND      g0326(.a(new_n342_), .b(new_n338_), .O(new_n343_));
  OR       g0327(.a(new_n343_), .b(new_n332_), .O(new_n344_));
  AND      g0328(.a(new_n204_), .b(i_2_0_13_0), .O(new_n345_));
  AND      g0329(.a(new_n345_), .b(new_n344_), .O(new_n346_));
  AND      g0330(.a(i_2_0_16_0), .b(i_2_0_13_0), .O(new_n347_));
  NAND     g0331(.a(new_n347_), .b(new_n23_), .O(new_n348_));
  OR       g0332(.a(new_n135_), .b(new_n177_), .O(new_n349_));
  OR       g0333(.a(new_n349_), .b(new_n70_), .O(new_n350_));
  OR       g0334(.a(new_n350_), .b(new_n348_), .O(new_n351_));
  OR       g0335(.a(new_n207_), .b(new_n137_), .O(new_n352_));
  OR       g0336(.a(new_n225_), .b(i_2_0_49_0), .O(new_n353_));
  OR       g0337(.a(new_n353_), .b(new_n352_), .O(new_n354_));
  NAND     g0338(.a(new_n354_), .b(new_n351_), .O(new_n355_));
  OR       g0339(.a(new_n355_), .b(new_n346_), .O(new_n356_));
  OR       g0340(.a(new_n356_), .b(new_n331_), .O(new_n357_));
  OR       g0341(.a(new_n357_), .b(new_n302_), .O(new_n358_));
  OR       g0342(.a(new_n358_), .b(new_n273_), .O(new_n359_));
  OR       g0343(.a(new_n359_), .b(new_n239_), .O(new_n360_));
  AND      g0344(.a(new_n360_), .b(new_n18_), .O(new_n361_));
  NOT      g0345(.a(i_2_0_66_0), .O(new_n362_));
  OR       g0346(.a(i_2_0_139_0), .b(new_n362_), .O(new_n363_));
  NOT      g0347(.a(new_n363_), .O(new_n364_));
  NAND     g0348(.a(new_n79_), .b(i_2_0_94_0), .O(new_n365_));
  OR       g0349(.a(new_n29_), .b(i_2_0_94_0), .O(new_n366_));
  OR       g0350(.a(new_n48_), .b(i_2_0_94_0), .O(new_n367_));
  NAND     g0351(.a(new_n367_), .b(new_n366_), .O(new_n368_));
  OR       g0352(.a(new_n368_), .b(new_n23_), .O(new_n369_));
  AND      g0353(.a(new_n369_), .b(new_n68_), .O(new_n370_));
  OR       g0354(.a(i_2_0_142_0), .b(i_2_0_94_0), .O(new_n371_));
  NOT      g0355(.a(new_n371_), .O(new_n372_));
  OR       g0356(.a(new_n372_), .b(new_n149_), .O(new_n373_));
  OR       g0357(.a(new_n25_), .b(new_n152_), .O(new_n374_));
  AND      g0358(.a(new_n374_), .b(new_n91_), .O(new_n375_));
  AND      g0359(.a(new_n375_), .b(new_n373_), .O(new_n376_));
  OR       g0360(.a(new_n376_), .b(new_n370_), .O(new_n377_));
  AND      g0361(.a(new_n377_), .b(new_n365_), .O(new_n378_));
  AND      g0362(.a(new_n82_), .b(i_2_0_13_0), .O(new_n379_));
  AND      g0363(.a(new_n48_), .b(new_n62_), .O(new_n380_));
  AND      g0364(.a(new_n380_), .b(new_n379_), .O(new_n381_));
  OR       g0365(.a(new_n381_), .b(new_n187_), .O(new_n382_));
  OR       g0366(.a(i_2_0_147_0), .b(i_2_0_94_0), .O(new_n383_));
  OR       g0367(.a(new_n383_), .b(new_n78_), .O(new_n384_));
  NAND     g0368(.a(i_2_0_109_0), .b(i_2_0_13_0), .O(new_n385_));
  AND      g0369(.a(new_n385_), .b(i_2_0_142_0), .O(new_n386_));
  NAND     g0370(.a(new_n386_), .b(new_n384_), .O(new_n387_));
  AND      g0371(.a(new_n387_), .b(new_n382_), .O(new_n388_));
  OR       g0372(.a(i_2_0_78_0), .b(new_n41_), .O(new_n389_));
  NOT      g0373(.a(new_n389_), .O(new_n390_));
  OR       g0374(.a(i_2_0_109_0), .b(i_2_0_94_0), .O(new_n391_));
  OR       g0375(.a(new_n391_), .b(new_n35_), .O(new_n392_));
  NAND     g0376(.a(new_n392_), .b(new_n105_), .O(new_n393_));
  AND      g0377(.a(new_n393_), .b(new_n390_), .O(new_n394_));
  AND      g0378(.a(new_n368_), .b(new_n229_), .O(new_n395_));
  OR       g0379(.a(new_n395_), .b(new_n394_), .O(new_n396_));
  OR       g0380(.a(new_n396_), .b(new_n388_), .O(new_n397_));
  OR       g0381(.a(new_n397_), .b(new_n378_), .O(new_n398_));
  AND      g0382(.a(new_n398_), .b(new_n364_), .O(new_n399_));
  AND      g0383(.a(new_n18_), .b(i_2_0_16_0), .O(new_n400_));
  NOT      g0384(.a(new_n137_), .O(new_n401_));
  AND      g0385(.a(i_2_0_109_0), .b(i_2_0_78_0), .O(new_n402_));
  OR       g0386(.a(new_n402_), .b(new_n401_), .O(new_n403_));
  NAND     g0387(.a(new_n403_), .b(new_n375_), .O(new_n404_));
  NAND     g0388(.a(new_n404_), .b(new_n241_), .O(new_n405_));
  AND      g0389(.a(new_n405_), .b(new_n400_), .O(new_n406_));
  OR       g0390(.a(i_2_0_139_0), .b(i_2_0_97_0), .O(new_n407_));
  OR       g0391(.a(new_n407_), .b(new_n51_), .O(new_n408_));
  OR       g0392(.a(new_n408_), .b(new_n29_), .O(new_n409_));
  NAND     g0393(.a(i_2_0_139_0), .b(i_2_0_97_0), .O(new_n410_));
  OR       g0394(.a(new_n410_), .b(new_n230_), .O(new_n411_));
  NAND     g0395(.a(new_n411_), .b(new_n368_), .O(new_n412_));
  NAND     g0396(.a(new_n412_), .b(new_n409_), .O(new_n413_));
  AND      g0397(.a(new_n413_), .b(new_n390_), .O(new_n414_));
  NAND     g0398(.a(new_n51_), .b(new_n71_), .O(new_n415_));
  OR       g0399(.a(new_n29_), .b(i_2_0_97_0), .O(new_n416_));
  NOT      g0400(.a(new_n416_), .O(new_n417_));
  OR       g0401(.a(i_2_0_94_0), .b(i_2_0_78_0), .O(new_n418_));
  NOT      g0402(.a(new_n418_), .O(new_n419_));
  AND      g0403(.a(new_n419_), .b(new_n417_), .O(new_n420_));
  AND      g0404(.a(new_n420_), .b(new_n415_), .O(new_n421_));
  OR       g0405(.a(new_n421_), .b(new_n414_), .O(new_n422_));
  OR       g0406(.a(new_n422_), .b(new_n406_), .O(new_n423_));
  AND      g0407(.a(new_n423_), .b(new_n82_), .O(new_n424_));
  OR       g0408(.a(new_n424_), .b(new_n399_), .O(new_n425_));
  OR       g0409(.a(new_n189_), .b(i_2_0_109_0), .O(new_n426_));
  NOT      g0410(.a(new_n426_), .O(new_n427_));
  NAND     g0411(.a(new_n224_), .b(i_2_0_94_0), .O(new_n428_));
  OR       g0412(.a(new_n428_), .b(new_n427_), .O(new_n429_));
  AND      g0413(.a(new_n429_), .b(new_n82_), .O(new_n430_));
  NOT      g0414(.a(new_n49_), .O(new_n431_));
  AND      g0415(.a(new_n431_), .b(new_n335_), .O(new_n432_));
  NAND     g0416(.a(new_n418_), .b(new_n383_), .O(new_n433_));
  NAND     g0417(.a(new_n19_), .b(new_n29_), .O(new_n434_));
  AND      g0418(.a(new_n434_), .b(new_n433_), .O(new_n435_));
  OR       g0419(.a(i_2_0_94_0), .b(new_n41_), .O(new_n436_));
  OR       g0420(.a(new_n436_), .b(i_2_0_109_0), .O(new_n437_));
  NAND     g0421(.a(new_n437_), .b(new_n389_), .O(new_n438_));
  OR       g0422(.a(new_n438_), .b(new_n435_), .O(new_n439_));
  OR       g0423(.a(new_n439_), .b(new_n432_), .O(new_n440_));
  OR       g0424(.a(new_n440_), .b(new_n430_), .O(new_n441_));
  AND      g0425(.a(new_n441_), .b(new_n364_), .O(new_n442_));
  AND      g0426(.a(i_2_0_147_0), .b(i_2_0_78_0), .O(new_n443_));
  OR       g0427(.a(new_n443_), .b(i_2_0_109_0), .O(new_n444_));
  AND      g0428(.a(new_n189_), .b(new_n29_), .O(new_n445_));
  AND      g0429(.a(new_n445_), .b(new_n444_), .O(new_n446_));
  NAND     g0430(.a(new_n372_), .b(new_n26_), .O(new_n447_));
  OR       g0431(.a(new_n447_), .b(new_n446_), .O(new_n448_));
  OR       g0432(.a(i_2_0_118_0), .b(new_n23_), .O(new_n449_));
  OR       g0433(.a(new_n449_), .b(new_n20_), .O(new_n450_));
  NAND     g0434(.a(new_n450_), .b(new_n372_), .O(new_n451_));
  AND      g0435(.a(new_n451_), .b(new_n41_), .O(new_n452_));
  NAND     g0436(.a(new_n419_), .b(new_n449_), .O(new_n453_));
  AND      g0437(.a(new_n453_), .b(i_2_0_142_0), .O(new_n454_));
  OR       g0438(.a(new_n372_), .b(new_n153_), .O(new_n455_));
  NAND     g0439(.a(new_n455_), .b(new_n21_), .O(new_n456_));
  OR       g0440(.a(new_n456_), .b(new_n454_), .O(new_n457_));
  OR       g0441(.a(new_n457_), .b(new_n452_), .O(new_n458_));
  NAND     g0442(.a(new_n458_), .b(new_n448_), .O(new_n459_));
  OR       g0443(.a(new_n228_), .b(new_n153_), .O(new_n460_));
  NAND     g0444(.a(i_2_0_109_0), .b(i_2_0_16_0), .O(new_n461_));
  AND      g0445(.a(new_n461_), .b(new_n371_), .O(new_n462_));
  OR       g0446(.a(new_n462_), .b(new_n402_), .O(new_n463_));
  NAND     g0447(.a(new_n463_), .b(new_n460_), .O(new_n464_));
  AND      g0448(.a(new_n464_), .b(new_n177_), .O(new_n465_));
  AND      g0449(.a(new_n20_), .b(new_n91_), .O(new_n466_));
  OR       g0450(.a(new_n466_), .b(new_n433_), .O(new_n467_));
  OR       g0451(.a(new_n25_), .b(new_n18_), .O(new_n468_));
  AND      g0452(.a(new_n468_), .b(new_n23_), .O(new_n469_));
  OR       g0453(.a(new_n469_), .b(new_n467_), .O(new_n470_));
  AND      g0454(.a(new_n470_), .b(new_n149_), .O(new_n471_));
  OR       g0455(.a(new_n471_), .b(new_n465_), .O(new_n472_));
  OR       g0456(.a(new_n472_), .b(new_n459_), .O(new_n473_));
  OR       g0457(.a(new_n473_), .b(new_n442_), .O(new_n474_));
  AND      g0458(.a(new_n474_), .b(i_2_0_13_0), .O(new_n475_));
  OR       g0459(.a(new_n475_), .b(new_n425_), .O(new_n476_));
  AND      g0460(.a(new_n33_), .b(i_2_0_66_0), .O(new_n477_));
  OR       g0461(.a(new_n371_), .b(i_2_0_109_0), .O(new_n478_));
  OR       g0462(.a(new_n45_), .b(new_n78_), .O(new_n479_));
  NAND     g0463(.a(new_n479_), .b(new_n478_), .O(new_n480_));
  OR       g0464(.a(new_n383_), .b(new_n29_), .O(new_n481_));
  AND      g0465(.a(new_n189_), .b(i_2_0_97_0), .O(new_n482_));
  NAND     g0466(.a(new_n482_), .b(new_n481_), .O(new_n483_));
  AND      g0467(.a(new_n483_), .b(new_n480_), .O(new_n484_));
  AND      g0468(.a(i_2_0_94_0), .b(new_n41_), .O(new_n485_));
  AND      g0469(.a(new_n485_), .b(new_n293_), .O(new_n486_));
  OR       g0470(.a(new_n170_), .b(new_n23_), .O(new_n487_));
  NAND     g0471(.a(new_n487_), .b(new_n264_), .O(new_n488_));
  OR       g0472(.a(new_n488_), .b(new_n486_), .O(new_n489_));
  AND      g0473(.a(new_n419_), .b(i_2_0_97_0), .O(new_n490_));
  NAND     g0474(.a(new_n490_), .b(new_n230_), .O(new_n491_));
  NAND     g0475(.a(new_n491_), .b(new_n489_), .O(new_n492_));
  OR       g0476(.a(i_2_0_139_0), .b(i_2_0_94_0), .O(new_n493_));
  NAND     g0477(.a(new_n493_), .b(new_n43_), .O(new_n494_));
  AND      g0478(.a(new_n494_), .b(new_n82_), .O(new_n495_));
  AND      g0479(.a(new_n229_), .b(new_n164_), .O(new_n496_));
  NAND     g0480(.a(new_n485_), .b(new_n277_), .O(new_n497_));
  AND      g0481(.a(new_n497_), .b(new_n496_), .O(new_n498_));
  OR       g0482(.a(new_n498_), .b(new_n495_), .O(new_n499_));
  OR       g0483(.a(new_n499_), .b(new_n492_), .O(new_n500_));
  OR       g0484(.a(new_n500_), .b(new_n484_), .O(new_n501_));
  OR       g0485(.a(new_n189_), .b(new_n21_), .O(new_n502_));
  OR       g0486(.a(i_2_0_118_0), .b(new_n63_), .O(new_n503_));
  OR       g0487(.a(i_2_0_97_0), .b(new_n18_), .O(new_n504_));
  OR       g0488(.a(new_n504_), .b(new_n503_), .O(new_n505_));
  NAND     g0489(.a(new_n505_), .b(new_n502_), .O(new_n506_));
  AND      g0490(.a(new_n506_), .b(new_n41_), .O(new_n507_));
  OR       g0491(.a(new_n443_), .b(new_n105_), .O(new_n508_));
  NAND     g0492(.a(new_n508_), .b(i_2_0_139_0), .O(new_n509_));
  OR       g0493(.a(i_2_0_118_0), .b(i_2_0_97_0), .O(new_n510_));
  AND      g0494(.a(new_n383_), .b(i_2_0_142_0), .O(new_n511_));
  NAND     g0495(.a(new_n511_), .b(new_n510_), .O(new_n512_));
  AND      g0496(.a(new_n512_), .b(new_n509_), .O(new_n513_));
  OR       g0497(.a(new_n513_), .b(new_n507_), .O(new_n514_));
  AND      g0498(.a(new_n514_), .b(new_n305_), .O(new_n515_));
  NOT      g0499(.a(new_n407_), .O(new_n516_));
  OR       g0500(.a(new_n279_), .b(new_n516_), .O(new_n517_));
  NAND     g0501(.a(new_n150_), .b(i_2_0_142_0), .O(new_n518_));
  AND      g0502(.a(new_n518_), .b(new_n517_), .O(new_n519_));
  OR       g0503(.a(new_n400_), .b(new_n373_), .O(new_n520_));
  NAND     g0504(.a(new_n253_), .b(i_2_0_78_0), .O(new_n521_));
  AND      g0505(.a(new_n521_), .b(new_n25_), .O(new_n522_));
  OR       g0506(.a(new_n522_), .b(new_n520_), .O(new_n523_));
  OR       g0507(.a(new_n523_), .b(new_n519_), .O(new_n524_));
  AND      g0508(.a(new_n524_), .b(i_2_0_13_0), .O(new_n525_));
  OR       g0509(.a(new_n525_), .b(new_n515_), .O(new_n526_));
  AND      g0510(.a(new_n152_), .b(i_2_0_16_0), .O(new_n527_));
  NAND     g0511(.a(new_n493_), .b(new_n28_), .O(new_n528_));
  AND      g0512(.a(new_n528_), .b(new_n164_), .O(new_n529_));
  OR       g0513(.a(new_n407_), .b(i_2_0_94_0), .O(new_n530_));
  OR       g0514(.a(new_n189_), .b(i_2_0_94_0), .O(new_n531_));
  NAND     g0515(.a(new_n531_), .b(new_n530_), .O(new_n532_));
  OR       g0516(.a(new_n532_), .b(new_n229_), .O(new_n533_));
  OR       g0517(.a(new_n533_), .b(new_n529_), .O(new_n534_));
  AND      g0518(.a(new_n534_), .b(new_n527_), .O(new_n535_));
  NAND     g0519(.a(i_2_0_97_0), .b(i_2_0_78_0), .O(new_n536_));
  NAND     g0520(.a(new_n436_), .b(new_n385_), .O(new_n537_));
  AND      g0521(.a(new_n537_), .b(new_n536_), .O(new_n538_));
  OR       g0522(.a(new_n496_), .b(new_n149_), .O(new_n539_));
  OR       g0523(.a(new_n539_), .b(new_n538_), .O(new_n540_));
  AND      g0524(.a(new_n540_), .b(new_n177_), .O(new_n541_));
  OR       g0525(.a(new_n541_), .b(new_n535_), .O(new_n542_));
  OR       g0526(.a(new_n542_), .b(new_n526_), .O(new_n543_));
  OR       g0527(.a(new_n543_), .b(new_n501_), .O(new_n544_));
  AND      g0528(.a(new_n544_), .b(new_n477_), .O(new_n545_));
  NOT      g0529(.a(new_n92_), .O(new_n546_));
  AND      g0530(.a(new_n365_), .b(i_2_0_66_0), .O(new_n547_));
  OR       g0531(.a(new_n78_), .b(i_2_0_139_0), .O(new_n548_));
  OR       g0532(.a(i_2_0_147_0), .b(new_n362_), .O(new_n549_));
  AND      g0533(.a(new_n549_), .b(new_n548_), .O(new_n550_));
  OR       g0534(.a(new_n261_), .b(i_2_0_97_0), .O(new_n551_));
  OR       g0535(.a(new_n551_), .b(new_n550_), .O(new_n552_));
  OR       g0536(.a(i_2_0_109_0), .b(new_n362_), .O(new_n553_));
  AND      g0537(.a(new_n553_), .b(i_2_0_94_0), .O(new_n554_));
  OR       g0538(.a(new_n554_), .b(i_2_0_139_0), .O(new_n555_));
  NAND     g0539(.a(new_n555_), .b(new_n552_), .O(new_n556_));
  OR       g0540(.a(new_n556_), .b(new_n547_), .O(new_n557_));
  AND      g0541(.a(new_n557_), .b(new_n68_), .O(new_n558_));
  NAND     g0542(.a(new_n61_), .b(i_2_0_66_0), .O(new_n559_));
  NAND     g0543(.a(new_n559_), .b(new_n256_), .O(new_n560_));
  AND      g0544(.a(new_n410_), .b(i_2_0_118_0), .O(new_n561_));
  AND      g0545(.a(new_n561_), .b(new_n560_), .O(new_n562_));
  OR       g0546(.a(new_n383_), .b(i_2_0_118_0), .O(new_n563_));
  OR       g0547(.a(new_n493_), .b(new_n29_), .O(new_n564_));
  NAND     g0548(.a(new_n564_), .b(new_n563_), .O(new_n565_));
  OR       g0549(.a(new_n565_), .b(new_n562_), .O(new_n566_));
  AND      g0550(.a(new_n566_), .b(new_n82_), .O(new_n567_));
  OR       g0551(.a(new_n416_), .b(new_n104_), .O(new_n568_));
  OR       g0552(.a(new_n51_), .b(new_n104_), .O(new_n569_));
  NAND     g0553(.a(new_n569_), .b(new_n568_), .O(new_n570_));
  OR       g0554(.a(new_n44_), .b(i_2_0_97_0), .O(new_n571_));
  OR       g0555(.a(i_2_0_97_0), .b(new_n362_), .O(new_n572_));
  OR       g0556(.a(new_n572_), .b(new_n391_), .O(new_n573_));
  NAND     g0557(.a(new_n573_), .b(new_n571_), .O(new_n574_));
  OR       g0558(.a(new_n574_), .b(new_n570_), .O(new_n575_));
  AND      g0559(.a(new_n575_), .b(new_n62_), .O(new_n576_));
  NOT      g0560(.a(new_n314_), .O(new_n577_));
  OR       g0561(.a(new_n35_), .b(new_n362_), .O(new_n578_));
  OR       g0562(.a(new_n253_), .b(i_2_0_16_0), .O(new_n579_));
  OR       g0563(.a(new_n579_), .b(new_n578_), .O(new_n580_));
  NAND     g0564(.a(new_n580_), .b(new_n478_), .O(new_n581_));
  AND      g0565(.a(new_n581_), .b(new_n577_), .O(new_n582_));
  OR       g0566(.a(new_n22_), .b(i_2_0_66_0), .O(new_n583_));
  OR       g0567(.a(new_n156_), .b(i_2_0_142_0), .O(new_n584_));
  NAND     g0568(.a(new_n584_), .b(new_n44_), .O(new_n585_));
  NAND     g0569(.a(new_n585_), .b(new_n583_), .O(new_n586_));
  NAND     g0570(.a(new_n586_), .b(new_n384_), .O(new_n587_));
  OR       g0571(.a(new_n587_), .b(new_n582_), .O(new_n588_));
  OR       g0572(.a(new_n588_), .b(new_n576_), .O(new_n589_));
  OR       g0573(.a(new_n589_), .b(new_n567_), .O(new_n590_));
  OR       g0574(.a(new_n590_), .b(new_n558_), .O(new_n591_));
  AND      g0575(.a(new_n591_), .b(new_n546_), .O(new_n592_));
  OR       g0576(.a(new_n592_), .b(new_n545_), .O(new_n593_));
  OR       g0577(.a(new_n593_), .b(new_n476_), .O(new_n594_));
  OR       g0578(.a(new_n285_), .b(i_2_0_16_0), .O(new_n595_));
  NAND     g0579(.a(i_2_0_109_0), .b(i_2_0_97_0), .O(new_n596_));
  AND      g0580(.a(new_n596_), .b(new_n24_), .O(new_n597_));
  AND      g0581(.a(new_n597_), .b(new_n595_), .O(new_n598_));
  OR       g0582(.a(i_2_0_16_0), .b(i_2_0_13_0), .O(new_n599_));
  AND      g0583(.a(new_n599_), .b(new_n289_), .O(new_n600_));
  NOT      g0584(.a(new_n347_), .O(new_n601_));
  OR       g0585(.a(new_n150_), .b(new_n78_), .O(new_n602_));
  NAND     g0586(.a(new_n602_), .b(new_n601_), .O(new_n603_));
  OR       g0587(.a(new_n603_), .b(new_n600_), .O(new_n604_));
  OR       g0588(.a(new_n604_), .b(new_n598_), .O(new_n605_));
  AND      g0589(.a(new_n605_), .b(new_n372_), .O(new_n606_));
  NAND     g0590(.a(new_n407_), .b(i_2_0_94_0), .O(new_n607_));
  NAND     g0591(.a(new_n607_), .b(new_n599_), .O(new_n608_));
  NAND     g0592(.a(new_n608_), .b(new_n530_), .O(new_n609_));
  AND      g0593(.a(new_n609_), .b(new_n111_), .O(new_n610_));
  OR       g0594(.a(new_n436_), .b(new_n228_), .O(new_n611_));
  NAND     g0595(.a(new_n347_), .b(new_n21_), .O(new_n612_));
  OR       g0596(.a(new_n612_), .b(new_n391_), .O(new_n613_));
  NAND     g0597(.a(new_n613_), .b(new_n611_), .O(new_n614_));
  OR       g0598(.a(new_n614_), .b(new_n610_), .O(new_n615_));
  AND      g0599(.a(new_n615_), .b(new_n164_), .O(new_n616_));
  AND      g0600(.a(new_n170_), .b(new_n21_), .O(new_n617_));
  OR       g0601(.a(new_n305_), .b(new_n617_), .O(new_n618_));
  NAND     g0602(.a(new_n612_), .b(new_n437_), .O(new_n619_));
  OR       g0603(.a(new_n619_), .b(new_n618_), .O(new_n620_));
  AND      g0604(.a(new_n373_), .b(new_n23_), .O(new_n621_));
  NAND     g0605(.a(new_n621_), .b(new_n620_), .O(new_n622_));
  OR       g0606(.a(new_n530_), .b(new_n601_), .O(new_n623_));
  NAND     g0607(.a(new_n623_), .b(new_n622_), .O(new_n624_));
  OR       g0608(.a(new_n624_), .b(new_n616_), .O(new_n625_));
  OR       g0609(.a(new_n625_), .b(new_n606_), .O(new_n626_));
  AND      g0610(.a(new_n626_), .b(new_n33_), .O(new_n627_));
  NAND     g0611(.a(new_n51_), .b(i_2_0_78_0), .O(new_n628_));
  AND      g0612(.a(new_n418_), .b(new_n41_), .O(new_n629_));
  NAND     g0613(.a(new_n629_), .b(new_n416_), .O(new_n630_));
  AND      g0614(.a(new_n630_), .b(new_n628_), .O(new_n631_));
  OR       g0615(.a(new_n485_), .b(i_2_0_97_0), .O(new_n632_));
  OR       g0616(.a(new_n51_), .b(new_n124_), .O(new_n633_));
  AND      g0617(.a(new_n633_), .b(new_n632_), .O(new_n634_));
  NAND     g0618(.a(new_n634_), .b(new_n367_), .O(new_n635_));
  OR       g0619(.a(new_n635_), .b(new_n631_), .O(new_n636_));
  AND      g0620(.a(new_n636_), .b(new_n379_), .O(new_n637_));
  NOT      g0621(.a(new_n383_), .O(new_n638_));
  AND      g0622(.a(new_n279_), .b(new_n211_), .O(new_n639_));
  OR       g0623(.a(new_n639_), .b(new_n638_), .O(new_n640_));
  AND      g0624(.a(new_n640_), .b(new_n347_), .O(new_n641_));
  OR       g0625(.a(new_n249_), .b(new_n23_), .O(new_n642_));
  AND      g0626(.a(new_n170_), .b(i_2_0_16_0), .O(new_n643_));
  AND      g0627(.a(new_n643_), .b(new_n18_), .O(new_n644_));
  AND      g0628(.a(new_n644_), .b(new_n642_), .O(new_n645_));
  OR       g0629(.a(new_n645_), .b(new_n641_), .O(new_n646_));
  OR       g0630(.a(new_n646_), .b(new_n637_), .O(new_n647_));
  NAND     g0631(.a(new_n531_), .b(new_n389_), .O(new_n648_));
  AND      g0632(.a(new_n648_), .b(new_n374_), .O(new_n649_));
  NAND     g0633(.a(new_n384_), .b(new_n224_), .O(new_n650_));
  AND      g0634(.a(new_n650_), .b(new_n649_), .O(new_n651_));
  OR       g0635(.a(new_n651_), .b(new_n400_), .O(new_n652_));
  AND      g0636(.a(new_n652_), .b(new_n82_), .O(new_n653_));
  OR       g0637(.a(new_n134_), .b(new_n18_), .O(new_n654_));
  AND      g0638(.a(new_n654_), .b(new_n230_), .O(new_n655_));
  OR       g0639(.a(new_n655_), .b(new_n649_), .O(new_n656_));
  AND      g0640(.a(new_n656_), .b(new_n229_), .O(new_n657_));
  OR       g0641(.a(new_n657_), .b(new_n653_), .O(new_n658_));
  OR       g0642(.a(new_n658_), .b(new_n647_), .O(new_n659_));
  AND      g0643(.a(new_n659_), .b(i_2_0_66_0), .O(new_n660_));
  OR       g0644(.a(i_2_0_147_0), .b(i_2_0_74_0), .O(new_n661_));
  NOT      g0645(.a(new_n661_), .O(new_n662_));
  NAND     g0646(.a(new_n548_), .b(new_n241_), .O(new_n663_));
  AND      g0647(.a(new_n663_), .b(new_n390_), .O(new_n664_));
  OR       g0648(.a(new_n255_), .b(new_n247_), .O(new_n665_));
  OR       g0649(.a(new_n632_), .b(new_n137_), .O(new_n666_));
  NAND     g0650(.a(new_n666_), .b(new_n665_), .O(new_n667_));
  OR       g0651(.a(new_n667_), .b(new_n664_), .O(new_n668_));
  AND      g0652(.a(new_n668_), .b(new_n82_), .O(new_n669_));
  OR       g0653(.a(new_n418_), .b(new_n410_), .O(new_n670_));
  OR       g0654(.a(new_n670_), .b(new_n247_), .O(new_n671_));
  NAND     g0655(.a(new_n671_), .b(new_n568_), .O(new_n672_));
  AND      g0656(.a(new_n672_), .b(i_2_0_57_0), .O(new_n673_));
  OR       g0657(.a(new_n126_), .b(i_2_0_118_0), .O(new_n674_));
  NAND     g0658(.a(new_n674_), .b(i_2_0_139_0), .O(new_n675_));
  AND      g0659(.a(new_n675_), .b(new_n379_), .O(new_n676_));
  NAND     g0660(.a(i_2_0_139_0), .b(i_2_0_16_0), .O(new_n677_));
  NAND     g0661(.a(new_n677_), .b(new_n42_), .O(new_n678_));
  AND      g0662(.a(new_n678_), .b(new_n490_), .O(new_n679_));
  OR       g0663(.a(new_n679_), .b(new_n676_), .O(new_n680_));
  OR       g0664(.a(new_n680_), .b(new_n673_), .O(new_n681_));
  AND      g0665(.a(new_n681_), .b(i_2_0_109_0), .O(new_n682_));
  AND      g0666(.a(new_n29_), .b(i_2_0_94_0), .O(new_n683_));
  AND      g0667(.a(new_n683_), .b(i_2_0_13_0), .O(new_n684_));
  OR       g0668(.a(new_n684_), .b(new_n643_), .O(new_n685_));
  AND      g0669(.a(new_n685_), .b(new_n516_), .O(new_n686_));
  OR       g0670(.a(new_n686_), .b(new_n682_), .O(new_n687_));
  OR       g0671(.a(new_n687_), .b(new_n669_), .O(new_n688_));
  AND      g0672(.a(new_n688_), .b(new_n662_), .O(new_n689_));
  OR       g0673(.a(new_n689_), .b(new_n660_), .O(new_n690_));
  OR       g0674(.a(new_n690_), .b(new_n627_), .O(new_n691_));
  OR       g0675(.a(new_n691_), .b(new_n594_), .O(new_n692_));
  AND      g0676(.a(new_n692_), .b(i_2_0_49_0), .O(new_n693_));
  AND      g0677(.a(new_n23_), .b(i_2_0_78_0), .O(new_n694_));
  AND      g0678(.a(new_n694_), .b(new_n230_), .O(new_n695_));
  NAND     g0679(.a(new_n551_), .b(new_n319_), .O(new_n696_));
  AND      g0680(.a(new_n696_), .b(new_n62_), .O(new_n697_));
  OR       g0681(.a(new_n697_), .b(new_n695_), .O(new_n698_));
  AND      g0682(.a(new_n698_), .b(new_n662_), .O(new_n699_));
  OR       g0683(.a(new_n314_), .b(new_n77_), .O(new_n700_));
  OR       g0684(.a(i_2_0_118_0), .b(i_2_0_109_0), .O(new_n701_));
  NAND     g0685(.a(new_n701_), .b(i_2_0_74_0), .O(new_n702_));
  NAND     g0686(.a(new_n702_), .b(new_n516_), .O(new_n703_));
  NAND     g0687(.a(new_n703_), .b(new_n700_), .O(new_n704_));
  OR       g0688(.a(new_n704_), .b(new_n699_), .O(new_n705_));
  AND      g0689(.a(new_n705_), .b(new_n64_), .O(new_n706_));
  OR       g0690(.a(new_n153_), .b(new_n124_), .O(new_n707_));
  NAND     g0691(.a(new_n707_), .b(new_n92_), .O(new_n708_));
  AND      g0692(.a(new_n708_), .b(new_n21_), .O(new_n709_));
  OR       g0693(.a(new_n154_), .b(i_2_0_74_0), .O(new_n710_));
  OR       g0694(.a(new_n710_), .b(new_n79_), .O(new_n711_));
  OR       g0695(.a(i_2_0_97_0), .b(i_2_0_57_0), .O(new_n712_));
  OR       g0696(.a(new_n712_), .b(new_n62_), .O(new_n713_));
  NAND     g0697(.a(new_n713_), .b(new_n711_), .O(new_n714_));
  OR       g0698(.a(new_n113_), .b(new_n152_), .O(new_n715_));
  NAND     g0699(.a(new_n715_), .b(new_n416_), .O(new_n716_));
  AND      g0700(.a(new_n716_), .b(new_n33_), .O(new_n717_));
  OR       g0701(.a(new_n717_), .b(new_n714_), .O(new_n718_));
  OR       g0702(.a(new_n718_), .b(new_n709_), .O(new_n719_));
  AND      g0703(.a(new_n336_), .b(i_2_0_97_0), .O(new_n720_));
  NAND     g0704(.a(i_2_0_118_0), .b(i_2_0_97_0), .O(new_n721_));
  NAND     g0705(.a(new_n721_), .b(new_n33_), .O(new_n722_));
  OR       g0706(.a(new_n722_), .b(new_n720_), .O(new_n723_));
  OR       g0707(.a(new_n218_), .b(new_n97_), .O(new_n724_));
  NAND     g0708(.a(new_n724_), .b(new_n723_), .O(new_n725_));
  AND      g0709(.a(new_n725_), .b(new_n401_), .O(new_n726_));
  OR       g0710(.a(new_n152_), .b(i_2_0_97_0), .O(new_n727_));
  AND      g0711(.a(new_n727_), .b(new_n79_), .O(new_n728_));
  NAND     g0712(.a(new_n311_), .b(new_n170_), .O(new_n729_));
  NAND     g0713(.a(new_n729_), .b(new_n728_), .O(new_n730_));
  AND      g0714(.a(new_n730_), .b(new_n63_), .O(new_n731_));
  OR       g0715(.a(new_n731_), .b(new_n726_), .O(new_n732_));
  OR       g0716(.a(new_n732_), .b(new_n719_), .O(new_n733_));
  AND      g0717(.a(new_n733_), .b(new_n347_), .O(new_n734_));
  NAND     g0718(.a(new_n164_), .b(i_2_0_109_0), .O(new_n735_));
  AND      g0719(.a(new_n735_), .b(new_n63_), .O(new_n736_));
  AND      g0720(.a(new_n170_), .b(i_2_0_147_0), .O(new_n737_));
  OR       g0721(.a(new_n737_), .b(new_n736_), .O(new_n738_));
  AND      g0722(.a(new_n738_), .b(new_n322_), .O(new_n739_));
  AND      g0723(.a(new_n739_), .b(new_n23_), .O(new_n740_));
  OR       g0724(.a(new_n740_), .b(new_n734_), .O(new_n741_));
  OR       g0725(.a(new_n741_), .b(new_n706_), .O(new_n742_));
  AND      g0726(.a(new_n742_), .b(new_n82_), .O(new_n743_));
  OR       g0727(.a(new_n715_), .b(new_n710_), .O(new_n744_));
  AND      g0728(.a(new_n205_), .b(new_n103_), .O(new_n745_));
  OR       g0729(.a(new_n97_), .b(i_2_0_78_0), .O(new_n746_));
  AND      g0730(.a(new_n746_), .b(new_n92_), .O(new_n747_));
  OR       g0731(.a(new_n747_), .b(new_n407_), .O(new_n748_));
  OR       g0732(.a(new_n748_), .b(new_n745_), .O(new_n749_));
  NAND     g0733(.a(new_n749_), .b(new_n744_), .O(new_n750_));
  AND      g0734(.a(new_n750_), .b(new_n347_), .O(new_n751_));
  OR       g0735(.a(new_n751_), .b(new_n743_), .O(new_n752_));
  NOT      g0736(.a(i_2_0_49_0), .O(new_n753_));
  OR       g0737(.a(i_2_0_57_0), .b(new_n753_), .O(new_n754_));
  NOT      g0738(.a(new_n754_), .O(new_n755_));
  AND      g0739(.a(new_n111_), .b(i_2_0_66_0), .O(new_n756_));
  OR       g0740(.a(new_n77_), .b(i_2_0_109_0), .O(new_n757_));
  OR       g0741(.a(new_n363_), .b(new_n152_), .O(new_n758_));
  NAND     g0742(.a(new_n758_), .b(new_n757_), .O(new_n759_));
  OR       g0743(.a(new_n759_), .b(new_n756_), .O(new_n760_));
  AND      g0744(.a(new_n760_), .b(new_n24_), .O(new_n761_));
  NOT      g0745(.a(new_n54_), .O(new_n762_));
  OR       g0746(.a(new_n153_), .b(i_2_0_147_0), .O(new_n763_));
  NAND     g0747(.a(new_n763_), .b(new_n551_), .O(new_n764_));
  AND      g0748(.a(new_n764_), .b(new_n762_), .O(new_n765_));
  OR       g0749(.a(i_2_0_142_0), .b(new_n362_), .O(new_n766_));
  OR       g0750(.a(new_n391_), .b(new_n77_), .O(new_n767_));
  NAND     g0751(.a(new_n767_), .b(new_n766_), .O(new_n768_));
  AND      g0752(.a(new_n768_), .b(new_n449_), .O(new_n769_));
  OR       g0753(.a(new_n510_), .b(new_n363_), .O(new_n770_));
  OR       g0754(.a(new_n42_), .b(i_2_0_142_0), .O(new_n771_));
  NAND     g0755(.a(new_n771_), .b(new_n770_), .O(new_n772_));
  OR       g0756(.a(new_n772_), .b(new_n769_), .O(new_n773_));
  OR       g0757(.a(new_n773_), .b(new_n765_), .O(new_n774_));
  OR       g0758(.a(new_n774_), .b(new_n761_), .O(new_n775_));
  AND      g0759(.a(new_n775_), .b(new_n62_), .O(new_n776_));
  OR       g0760(.a(new_n428_), .b(new_n69_), .O(new_n777_));
  OR       g0761(.a(i_2_0_94_0), .b(i_2_0_74_0), .O(new_n778_));
  NOT      g0762(.a(new_n778_), .O(new_n779_));
  NAND     g0763(.a(new_n391_), .b(new_n362_), .O(new_n780_));
  OR       g0764(.a(new_n780_), .b(new_n779_), .O(new_n781_));
  NAND     g0765(.a(new_n781_), .b(new_n777_), .O(new_n782_));
  NAND     g0766(.a(new_n782_), .b(new_n79_), .O(new_n783_));
  AND      g0767(.a(new_n783_), .b(new_n82_), .O(new_n784_));
  OR       g0768(.a(new_n78_), .b(i_2_0_142_0), .O(new_n785_));
  NAND     g0769(.a(new_n578_), .b(new_n785_), .O(new_n786_));
  AND      g0770(.a(new_n786_), .b(i_2_0_78_0), .O(new_n787_));
  OR       g0771(.a(new_n372_), .b(new_n22_), .O(new_n788_));
  AND      g0772(.a(new_n788_), .b(new_n23_), .O(new_n789_));
  NOT      g0773(.a(new_n493_), .O(new_n790_));
  AND      g0774(.a(new_n477_), .b(new_n790_), .O(new_n791_));
  AND      g0775(.a(new_n780_), .b(i_2_0_16_0), .O(new_n792_));
  OR       g0776(.a(new_n792_), .b(new_n791_), .O(new_n793_));
  OR       g0777(.a(new_n793_), .b(new_n789_), .O(new_n794_));
  OR       g0778(.a(new_n794_), .b(new_n787_), .O(new_n795_));
  OR       g0779(.a(new_n795_), .b(new_n784_), .O(new_n796_));
  OR       g0780(.a(new_n796_), .b(new_n776_), .O(new_n797_));
  AND      g0781(.a(new_n797_), .b(i_2_0_13_0), .O(new_n798_));
  OR       g0782(.a(new_n572_), .b(new_n485_), .O(new_n799_));
  NAND     g0783(.a(new_n799_), .b(new_n407_), .O(new_n800_));
  OR       g0784(.a(new_n780_), .b(i_2_0_16_0), .O(new_n801_));
  AND      g0785(.a(new_n801_), .b(new_n800_), .O(new_n802_));
  AND      g0786(.a(i_2_0_118_0), .b(i_2_0_66_0), .O(new_n803_));
  NAND     g0787(.a(new_n803_), .b(i_2_0_16_0), .O(new_n804_));
  NAND     g0788(.a(new_n804_), .b(new_n493_), .O(new_n805_));
  AND      g0789(.a(new_n805_), .b(new_n333_), .O(new_n806_));
  NAND     g0790(.a(new_n548_), .b(i_2_0_94_0), .O(new_n807_));
  AND      g0791(.a(new_n123_), .b(i_2_0_66_0), .O(new_n808_));
  AND      g0792(.a(new_n808_), .b(new_n807_), .O(new_n809_));
  OR       g0793(.a(new_n809_), .b(new_n806_), .O(new_n810_));
  OR       g0794(.a(new_n810_), .b(new_n802_), .O(new_n811_));
  AND      g0795(.a(new_n811_), .b(new_n82_), .O(new_n812_));
  OR       g0796(.a(new_n420_), .b(new_n400_), .O(new_n813_));
  AND      g0797(.a(new_n813_), .b(new_n364_), .O(new_n814_));
  OR       g0798(.a(new_n371_), .b(new_n211_), .O(new_n815_));
  OR       g0799(.a(new_n553_), .b(new_n293_), .O(new_n816_));
  NAND     g0800(.a(new_n816_), .b(new_n815_), .O(new_n817_));
  AND      g0801(.a(new_n817_), .b(i_2_0_74_0), .O(new_n818_));
  AND      g0802(.a(new_n695_), .b(i_2_0_66_0), .O(new_n819_));
  OR       g0803(.a(new_n819_), .b(new_n818_), .O(new_n820_));
  OR       g0804(.a(new_n820_), .b(new_n814_), .O(new_n821_));
  OR       g0805(.a(new_n821_), .b(new_n812_), .O(new_n822_));
  OR       g0806(.a(new_n822_), .b(new_n798_), .O(new_n823_));
  AND      g0807(.a(new_n823_), .b(new_n755_), .O(new_n824_));
  AND      g0808(.a(new_n516_), .b(new_n230_), .O(new_n825_));
  NOT      g0809(.a(new_n825_), .O(new_n826_));
  AND      g0810(.a(new_n551_), .b(i_2_0_78_0), .O(new_n827_));
  AND      g0811(.a(i_2_0_139_0), .b(new_n23_), .O(new_n828_));
  OR       g0812(.a(new_n828_), .b(new_n80_), .O(new_n829_));
  OR       g0813(.a(new_n829_), .b(new_n827_), .O(new_n830_));
  AND      g0814(.a(new_n830_), .b(new_n826_), .O(new_n831_));
  OR       g0815(.a(new_n831_), .b(i_2_0_74_0), .O(new_n832_));
  OR       g0816(.a(new_n261_), .b(new_n712_), .O(new_n833_));
  AND      g0817(.a(new_n833_), .b(new_n92_), .O(new_n834_));
  OR       g0818(.a(new_n97_), .b(i_2_0_139_0), .O(new_n835_));
  AND      g0819(.a(new_n835_), .b(new_n407_), .O(new_n836_));
  OR       g0820(.a(new_n836_), .b(new_n834_), .O(new_n837_));
  OR       g0821(.a(new_n30_), .b(new_n156_), .O(new_n838_));
  AND      g0822(.a(new_n757_), .b(new_n208_), .O(new_n839_));
  AND      g0823(.a(new_n839_), .b(new_n838_), .O(new_n840_));
  OR       g0824(.a(new_n840_), .b(new_n75_), .O(new_n841_));
  OR       g0825(.a(new_n255_), .b(new_n137_), .O(new_n842_));
  AND      g0826(.a(new_n156_), .b(i_2_0_97_0), .O(new_n843_));
  OR       g0827(.a(new_n843_), .b(new_n19_), .O(new_n844_));
  OR       g0828(.a(new_n844_), .b(new_n138_), .O(new_n845_));
  AND      g0829(.a(new_n845_), .b(new_n842_), .O(new_n846_));
  AND      g0830(.a(new_n846_), .b(new_n841_), .O(new_n847_));
  AND      g0831(.a(new_n847_), .b(new_n837_), .O(new_n848_));
  NAND     g0832(.a(new_n848_), .b(new_n832_), .O(new_n849_));
  AND      g0833(.a(new_n849_), .b(new_n379_), .O(new_n850_));
  OR       g0834(.a(new_n628_), .b(new_n516_), .O(new_n851_));
  AND      g0835(.a(new_n851_), .b(new_n561_), .O(new_n852_));
  NOT      g0836(.a(new_n91_), .O(new_n853_));
  AND      g0837(.a(i_2_0_109_0), .b(new_n62_), .O(new_n854_));
  OR       g0838(.a(new_n854_), .b(new_n260_), .O(new_n855_));
  AND      g0839(.a(new_n855_), .b(new_n853_), .O(new_n856_));
  NAND     g0840(.a(new_n35_), .b(i_2_0_57_0), .O(new_n857_));
  NAND     g0841(.a(new_n19_), .b(i_2_0_139_0), .O(new_n858_));
  AND      g0842(.a(new_n858_), .b(new_n857_), .O(new_n859_));
  AND      g0843(.a(new_n536_), .b(new_n401_), .O(new_n860_));
  OR       g0844(.a(new_n860_), .b(new_n859_), .O(new_n861_));
  OR       g0845(.a(new_n861_), .b(new_n856_), .O(new_n862_));
  OR       g0846(.a(new_n862_), .b(new_n852_), .O(new_n863_));
  AND      g0847(.a(new_n863_), .b(new_n149_), .O(new_n864_));
  NAND     g0848(.a(new_n228_), .b(new_n63_), .O(new_n865_));
  OR       g0849(.a(new_n596_), .b(i_2_0_147_0), .O(new_n866_));
  OR       g0850(.a(new_n866_), .b(new_n150_), .O(new_n867_));
  OR       g0851(.a(new_n720_), .b(i_2_0_142_0), .O(new_n868_));
  NAND     g0852(.a(new_n868_), .b(new_n867_), .O(new_n869_));
  AND      g0853(.a(new_n869_), .b(new_n865_), .O(new_n870_));
  NAND     g0854(.a(new_n426_), .b(new_n29_), .O(new_n871_));
  AND      g0855(.a(new_n871_), .b(new_n68_), .O(new_n872_));
  NOT      g0856(.a(new_n504_), .O(new_n873_));
  AND      g0857(.a(new_n873_), .b(new_n380_), .O(new_n874_));
  OR       g0858(.a(new_n874_), .b(new_n872_), .O(new_n875_));
  OR       g0859(.a(new_n875_), .b(new_n870_), .O(new_n876_));
  AND      g0860(.a(new_n876_), .b(new_n34_), .O(new_n877_));
  OR       g0861(.a(new_n877_), .b(new_n864_), .O(new_n878_));
  AND      g0862(.a(new_n878_), .b(i_2_0_13_0), .O(new_n879_));
  AND      g0863(.a(new_n838_), .b(i_2_0_57_0), .O(new_n880_));
  OR       g0864(.a(new_n880_), .b(new_n844_), .O(new_n881_));
  OR       g0865(.a(new_n24_), .b(i_2_0_74_0), .O(new_n882_));
  OR       g0866(.a(new_n882_), .b(new_n596_), .O(new_n883_));
  AND      g0867(.a(new_n35_), .b(new_n92_), .O(new_n884_));
  AND      g0868(.a(new_n884_), .b(new_n883_), .O(new_n885_));
  OR       g0869(.a(new_n885_), .b(new_n96_), .O(new_n886_));
  NAND     g0870(.a(new_n886_), .b(new_n881_), .O(new_n887_));
  AND      g0871(.a(new_n887_), .b(i_2_0_118_0), .O(new_n888_));
  OR       g0872(.a(new_n255_), .b(new_n77_), .O(new_n889_));
  AND      g0873(.a(new_n661_), .b(new_n75_), .O(new_n890_));
  OR       g0874(.a(new_n402_), .b(new_n407_), .O(new_n891_));
  OR       g0875(.a(new_n891_), .b(new_n890_), .O(new_n892_));
  NAND     g0876(.a(new_n892_), .b(new_n889_), .O(new_n893_));
  OR       g0877(.a(new_n893_), .b(new_n888_), .O(new_n894_));
  AND      g0878(.a(new_n894_), .b(new_n149_), .O(new_n895_));
  OR       g0879(.a(new_n895_), .b(new_n879_), .O(new_n896_));
  OR       g0880(.a(new_n896_), .b(new_n850_), .O(new_n897_));
  AND      g0881(.a(new_n897_), .b(i_2_0_66_0), .O(new_n898_));
  OR       g0882(.a(new_n898_), .b(new_n824_), .O(new_n899_));
  OR       g0883(.a(new_n899_), .b(new_n752_), .O(new_n900_));
  OR       g0884(.a(new_n900_), .b(new_n693_), .O(new_n901_));
  OR       g0885(.a(new_n901_), .b(new_n361_), .O(new_n902_));
  AND      g0886(.a(new_n902_), .b(new_n17_), .O(new_n903_));
  AND      g0887(.a(new_n756_), .b(new_n487_), .O(new_n904_));
  OR       g0888(.a(new_n175_), .b(new_n124_), .O(new_n905_));
  NAND     g0889(.a(new_n905_), .b(new_n28_), .O(new_n906_));
  NOT      g0890(.a(new_n766_), .O(new_n907_));
  XOR      g0891(.a(i_2_0_118_0), .b(i_2_0_109_0), .O(new_n908_));
  OR       g0892(.a(new_n908_), .b(new_n62_), .O(new_n909_));
  AND      g0893(.a(new_n909_), .b(new_n907_), .O(new_n910_));
  AND      g0894(.a(new_n496_), .b(i_2_0_109_0), .O(new_n911_));
  OR       g0895(.a(new_n911_), .b(new_n63_), .O(new_n912_));
  OR       g0896(.a(new_n912_), .b(new_n910_), .O(new_n913_));
  AND      g0897(.a(new_n913_), .b(new_n906_), .O(new_n914_));
  OR       g0898(.a(new_n914_), .b(new_n904_), .O(new_n915_));
  AND      g0899(.a(new_n915_), .b(new_n33_), .O(new_n916_));
  AND      g0900(.a(new_n907_), .b(new_n158_), .O(new_n917_));
  OR       g0901(.a(new_n150_), .b(new_n79_), .O(new_n918_));
  OR       g0902(.a(new_n918_), .b(i_2_0_142_0), .O(new_n919_));
  NAND     g0903(.a(new_n919_), .b(new_n191_), .O(new_n920_));
  OR       g0904(.a(new_n920_), .b(new_n917_), .O(new_n921_));
  AND      g0905(.a(new_n921_), .b(new_n23_), .O(new_n922_));
  NOT      g0906(.a(new_n138_), .O(new_n923_));
  NOT      g0907(.a(new_n553_), .O(new_n924_));
  OR       g0908(.a(new_n924_), .b(new_n854_), .O(new_n925_));
  AND      g0909(.a(new_n925_), .b(new_n923_), .O(new_n926_));
  NAND     g0910(.a(new_n858_), .b(new_n319_), .O(new_n927_));
  OR       g0911(.a(new_n927_), .b(new_n113_), .O(new_n928_));
  NAND     g0912(.a(new_n803_), .b(new_n628_), .O(new_n929_));
  OR       g0913(.a(new_n929_), .b(i_2_0_139_0), .O(new_n930_));
  NAND     g0914(.a(new_n930_), .b(new_n928_), .O(new_n931_));
  OR       g0915(.a(new_n931_), .b(new_n926_), .O(new_n932_));
  AND      g0916(.a(new_n932_), .b(new_n82_), .O(new_n933_));
  OR       g0917(.a(new_n933_), .b(new_n922_), .O(new_n934_));
  OR       g0918(.a(new_n934_), .b(new_n916_), .O(new_n935_));
  AND      g0919(.a(new_n935_), .b(i_2_0_49_0), .O(new_n936_));
  AND      g0920(.a(new_n83_), .b(new_n753_), .O(new_n937_));
  OR       g0921(.a(new_n402_), .b(new_n228_), .O(new_n938_));
  OR       g0922(.a(new_n938_), .b(new_n937_), .O(new_n939_));
  OR       g0923(.a(new_n720_), .b(new_n766_), .O(new_n940_));
  NAND     g0924(.a(new_n940_), .b(new_n939_), .O(new_n941_));
  NAND     g0925(.a(i_2_0_66_0), .b(i_2_0_49_0), .O(new_n942_));
  OR       g0926(.a(new_n942_), .b(new_n633_), .O(new_n943_));
  OR       g0927(.a(new_n754_), .b(new_n124_), .O(new_n944_));
  NAND     g0928(.a(new_n944_), .b(new_n943_), .O(new_n945_));
  OR       g0929(.a(new_n945_), .b(new_n941_), .O(new_n946_));
  AND      g0930(.a(new_n946_), .b(i_2_0_118_0), .O(new_n947_));
  OR       g0931(.a(i_2_0_109_0), .b(i_2_0_57_0), .O(new_n948_));
  OR       g0932(.a(new_n948_), .b(new_n753_), .O(new_n949_));
  OR       g0933(.a(new_n443_), .b(i_2_0_97_0), .O(new_n950_));
  OR       g0934(.a(new_n950_), .b(new_n949_), .O(new_n951_));
  NAND     g0935(.a(new_n951_), .b(new_n228_), .O(new_n952_));
  NAND     g0936(.a(new_n766_), .b(new_n444_), .O(new_n953_));
  AND      g0937(.a(new_n953_), .b(i_2_0_49_0), .O(new_n954_));
  OR       g0938(.a(new_n549_), .b(new_n402_), .O(new_n955_));
  NAND     g0939(.a(new_n955_), .b(i_2_0_57_0), .O(new_n956_));
  OR       g0940(.a(new_n956_), .b(new_n954_), .O(new_n957_));
  AND      g0941(.a(new_n957_), .b(new_n952_), .O(new_n958_));
  OR       g0942(.a(new_n958_), .b(new_n947_), .O(new_n959_));
  OR       g0943(.a(new_n948_), .b(new_n23_), .O(new_n960_));
  NAND     g0944(.a(new_n960_), .b(new_n67_), .O(new_n961_));
  AND      g0945(.a(new_n961_), .b(i_2_0_66_0), .O(new_n962_));
  OR       g0946(.a(i_2_0_57_0), .b(i_2_0_49_0), .O(new_n963_));
  NAND     g0947(.a(i_2_0_143_0), .b(i_2_0_78_0), .O(new_n964_));
  OR       g0948(.a(new_n964_), .b(new_n963_), .O(new_n965_));
  AND      g0949(.a(new_n596_), .b(new_n753_), .O(new_n966_));
  AND      g0950(.a(i_2_0_109_0), .b(i_2_0_49_0), .O(new_n967_));
  OR       g0951(.a(new_n967_), .b(new_n67_), .O(new_n968_));
  OR       g0952(.a(new_n968_), .b(new_n966_), .O(new_n969_));
  NAND     g0953(.a(new_n969_), .b(new_n965_), .O(new_n970_));
  OR       g0954(.a(new_n970_), .b(new_n962_), .O(new_n971_));
  AND      g0955(.a(new_n971_), .b(new_n25_), .O(new_n972_));
  OR       g0956(.a(new_n942_), .b(new_n28_), .O(new_n973_));
  OR       g0957(.a(new_n67_), .b(i_2_0_57_0), .O(new_n974_));
  NAND     g0958(.a(new_n974_), .b(new_n973_), .O(new_n975_));
  OR       g0959(.a(new_n975_), .b(new_n972_), .O(new_n976_));
  OR       g0960(.a(new_n976_), .b(new_n959_), .O(new_n977_));
  AND      g0961(.a(new_n977_), .b(new_n321_), .O(new_n978_));
  NAND     g0962(.a(new_n663_), .b(new_n62_), .O(new_n979_));
  NAND     g0963(.a(new_n979_), .b(new_n408_), .O(new_n980_));
  NOT      g0964(.a(new_n843_), .O(new_n981_));
  AND      g0965(.a(new_n981_), .b(new_n303_), .O(new_n982_));
  AND      g0966(.a(new_n982_), .b(new_n980_), .O(new_n983_));
  NAND     g0967(.a(new_n553_), .b(new_n416_), .O(new_n984_));
  AND      g0968(.a(new_n984_), .b(new_n76_), .O(new_n985_));
  OR       g0969(.a(i_2_0_109_0), .b(i_2_0_97_0), .O(new_n986_));
  OR       g0970(.a(new_n729_), .b(new_n986_), .O(new_n987_));
  OR       g0971(.a(new_n572_), .b(new_n224_), .O(new_n988_));
  NAND     g0972(.a(new_n988_), .b(new_n987_), .O(new_n989_));
  OR       g0973(.a(new_n989_), .b(new_n985_), .O(new_n990_));
  AND      g0974(.a(new_n990_), .b(new_n762_), .O(new_n991_));
  AND      g0975(.a(new_n62_), .b(i_2_0_66_0), .O(new_n992_));
  AND      g0976(.a(new_n992_), .b(new_n264_), .O(new_n993_));
  AND      g0977(.a(new_n993_), .b(new_n825_), .O(new_n994_));
  OR       g0978(.a(new_n994_), .b(new_n991_), .O(new_n995_));
  OR       g0979(.a(new_n995_), .b(new_n983_), .O(new_n996_));
  OR       g0980(.a(new_n996_), .b(new_n978_), .O(new_n997_));
  OR       g0981(.a(new_n997_), .b(new_n936_), .O(new_n998_));
  AND      g0982(.a(new_n998_), .b(new_n400_), .O(new_n999_));
  AND      g0983(.a(new_n321_), .b(i_2_0_66_0), .O(new_n1000_));
  AND      g0984(.a(new_n1000_), .b(new_n375_), .O(new_n1001_));
  OR       g0985(.a(new_n113_), .b(new_n29_), .O(new_n1002_));
  OR       g0986(.a(i_2_0_139_0), .b(i_2_0_57_0), .O(new_n1003_));
  AND      g0987(.a(new_n553_), .b(new_n661_), .O(new_n1004_));
  OR       g0988(.a(new_n1004_), .b(new_n1003_), .O(new_n1005_));
  NAND     g0989(.a(new_n1005_), .b(new_n1002_), .O(new_n1006_));
  OR       g0990(.a(new_n1006_), .b(new_n1001_), .O(new_n1007_));
  AND      g0991(.a(new_n1007_), .b(new_n23_), .O(new_n1008_));
  NOT      g0992(.a(new_n477_), .O(new_n1009_));
  OR       g0993(.a(new_n918_), .b(new_n1009_), .O(new_n1010_));
  OR       g0994(.a(new_n98_), .b(i_2_0_74_0), .O(new_n1011_));
  NAND     g0995(.a(new_n1011_), .b(new_n835_), .O(new_n1012_));
  AND      g0996(.a(new_n1012_), .b(new_n924_), .O(new_n1013_));
  OR       g0997(.a(new_n477_), .b(new_n63_), .O(new_n1014_));
  AND      g0998(.a(new_n1014_), .b(new_n349_), .O(new_n1015_));
  OR       g0999(.a(new_n1015_), .b(new_n1013_), .O(new_n1016_));
  NAND     g1000(.a(new_n1016_), .b(new_n132_), .O(new_n1017_));
  NAND     g1001(.a(new_n1017_), .b(new_n1010_), .O(new_n1018_));
  OR       g1002(.a(new_n1018_), .b(new_n1008_), .O(new_n1019_));
  AND      g1003(.a(new_n1019_), .b(i_2_0_49_0), .O(new_n1020_));
  OR       g1004(.a(new_n661_), .b(new_n120_), .O(new_n1021_));
  NAND     g1005(.a(new_n415_), .b(new_n33_), .O(new_n1022_));
  NAND     g1006(.a(new_n1022_), .b(new_n835_), .O(new_n1023_));
  NAND     g1007(.a(new_n1023_), .b(new_n992_), .O(new_n1024_));
  NAND     g1008(.a(new_n1024_), .b(new_n1021_), .O(new_n1025_));
  AND      g1009(.a(new_n1025_), .b(new_n755_), .O(new_n1026_));
  OR       g1010(.a(i_2_0_109_0), .b(i_2_0_74_0), .O(new_n1027_));
  OR       g1011(.a(new_n156_), .b(new_n362_), .O(new_n1028_));
  NAND     g1012(.a(new_n1028_), .b(new_n1027_), .O(new_n1029_));
  AND      g1013(.a(new_n1029_), .b(new_n694_), .O(new_n1030_));
  NOT      g1014(.a(new_n402_), .O(new_n1031_));
  AND      g1015(.a(new_n1031_), .b(i_2_0_147_0), .O(new_n1032_));
  AND      g1016(.a(new_n1032_), .b(new_n1000_), .O(new_n1033_));
  OR       g1017(.a(new_n1033_), .b(new_n1030_), .O(new_n1034_));
  AND      g1018(.a(new_n1034_), .b(new_n923_), .O(new_n1035_));
  OR       g1019(.a(new_n1035_), .b(new_n1026_), .O(new_n1036_));
  OR       g1020(.a(new_n1036_), .b(new_n1020_), .O(new_n1037_));
  AND      g1021(.a(new_n1037_), .b(new_n372_), .O(new_n1038_));
  AND      g1022(.a(new_n21_), .b(i_2_0_49_0), .O(new_n1039_));
  NOT      g1023(.a(new_n1027_), .O(new_n1040_));
  AND      g1024(.a(new_n536_), .b(new_n25_), .O(new_n1041_));
  NAND     g1025(.a(new_n124_), .b(new_n91_), .O(new_n1042_));
  OR       g1026(.a(new_n1042_), .b(new_n1041_), .O(new_n1043_));
  AND      g1027(.a(new_n1043_), .b(new_n1040_), .O(new_n1044_));
  NAND     g1028(.a(new_n211_), .b(new_n712_), .O(new_n1045_));
  AND      g1029(.a(new_n857_), .b(new_n33_), .O(new_n1046_));
  AND      g1030(.a(new_n1046_), .b(new_n1045_), .O(new_n1047_));
  AND      g1031(.a(new_n427_), .b(new_n31_), .O(new_n1048_));
  OR       g1032(.a(new_n1048_), .b(new_n1047_), .O(new_n1049_));
  OR       g1033(.a(new_n1049_), .b(new_n1044_), .O(new_n1050_));
  AND      g1034(.a(new_n1050_), .b(new_n1039_), .O(new_n1051_));
  OR       g1035(.a(new_n92_), .b(new_n23_), .O(new_n1052_));
  OR       g1036(.a(new_n754_), .b(i_2_0_78_0), .O(new_n1053_));
  OR       g1037(.a(new_n882_), .b(new_n124_), .O(new_n1054_));
  AND      g1038(.a(new_n1054_), .b(new_n1053_), .O(new_n1055_));
  NAND     g1039(.a(new_n1055_), .b(new_n1052_), .O(new_n1056_));
  AND      g1040(.a(new_n1056_), .b(new_n401_), .O(new_n1057_));
  AND      g1041(.a(i_2_0_118_0), .b(i_2_0_49_0), .O(new_n1058_));
  AND      g1042(.a(new_n1058_), .b(new_n63_), .O(new_n1059_));
  AND      g1043(.a(new_n340_), .b(new_n304_), .O(new_n1060_));
  AND      g1044(.a(new_n1060_), .b(new_n1059_), .O(new_n1061_));
  OR       g1045(.a(new_n1061_), .b(new_n1057_), .O(new_n1062_));
  OR       g1046(.a(new_n1062_), .b(new_n1051_), .O(new_n1063_));
  AND      g1047(.a(new_n1063_), .b(i_2_0_66_0), .O(new_n1064_));
  AND      g1048(.a(new_n153_), .b(new_n23_), .O(new_n1065_));
  NAND     g1049(.a(new_n1065_), .b(new_n171_), .O(new_n1066_));
  OR       g1050(.a(new_n1066_), .b(new_n927_), .O(new_n1067_));
  OR       g1051(.a(new_n248_), .b(i_2_0_139_0), .O(new_n1068_));
  NAND     g1052(.a(new_n1068_), .b(new_n1067_), .O(new_n1069_));
  AND      g1053(.a(new_n114_), .b(i_2_0_49_0), .O(new_n1070_));
  AND      g1054(.a(new_n1070_), .b(new_n1069_), .O(new_n1071_));
  OR       g1055(.a(new_n1071_), .b(new_n1064_), .O(new_n1072_));
  AND      g1056(.a(new_n1072_), .b(new_n149_), .O(new_n1073_));
  OR       g1057(.a(i_2_0_118_0), .b(new_n753_), .O(new_n1074_));
  OR       g1058(.a(new_n1074_), .b(new_n536_), .O(new_n1075_));
  NAND     g1059(.a(new_n1075_), .b(new_n255_), .O(new_n1076_));
  OR       g1060(.a(new_n77_), .b(i_2_0_142_0), .O(new_n1077_));
  NOT      g1061(.a(new_n1077_), .O(new_n1078_));
  OR       g1062(.a(new_n553_), .b(new_n113_), .O(new_n1079_));
  NOT      g1063(.a(new_n1079_), .O(new_n1080_));
  AND      g1064(.a(new_n1080_), .b(new_n1078_), .O(new_n1081_));
  AND      g1065(.a(new_n1081_), .b(new_n1076_), .O(new_n1082_));
  OR       g1066(.a(new_n1082_), .b(new_n1073_), .O(new_n1083_));
  OR       g1067(.a(new_n1083_), .b(new_n1038_), .O(new_n1084_));
  OR       g1068(.a(new_n1084_), .b(new_n999_), .O(new_n1085_));
  NAND     g1069(.a(new_n701_), .b(i_2_0_78_0), .O(new_n1086_));
  AND      g1070(.a(new_n1086_), .b(i_2_0_97_0), .O(new_n1087_));
  OR       g1071(.a(new_n1087_), .b(new_n135_), .O(new_n1088_));
  AND      g1072(.a(new_n1088_), .b(new_n33_), .O(new_n1089_));
  NOT      g1073(.a(new_n1058_), .O(new_n1090_));
  OR       g1074(.a(new_n1090_), .b(new_n51_), .O(new_n1091_));
  NAND     g1075(.a(new_n1091_), .b(new_n882_), .O(new_n1092_));
  OR       g1076(.a(new_n1092_), .b(new_n1089_), .O(new_n1093_));
  AND      g1077(.a(new_n1093_), .b(i_2_0_66_0), .O(new_n1094_));
  NAND     g1078(.a(new_n683_), .b(new_n854_), .O(new_n1095_));
  NAND     g1079(.a(new_n1095_), .b(new_n391_), .O(new_n1096_));
  OR       g1080(.a(new_n79_), .b(new_n168_), .O(new_n1097_));
  NAND     g1081(.a(new_n1097_), .b(new_n763_), .O(new_n1098_));
  OR       g1082(.a(new_n1098_), .b(new_n1096_), .O(new_n1099_));
  AND      g1083(.a(new_n1099_), .b(i_2_0_49_0), .O(new_n1100_));
  NOT      g1084(.a(new_n366_), .O(new_n1101_));
  AND      g1085(.a(new_n925_), .b(new_n1101_), .O(new_n1102_));
  OR       g1086(.a(new_n1102_), .b(new_n755_), .O(new_n1103_));
  NOT      g1087(.a(new_n180_), .O(new_n1104_));
  AND      g1088(.a(new_n1104_), .b(new_n230_), .O(new_n1105_));
  AND      g1089(.a(i_2_0_109_0), .b(new_n33_), .O(new_n1106_));
  OR       g1090(.a(new_n1106_), .b(new_n63_), .O(new_n1107_));
  AND      g1091(.a(new_n1107_), .b(new_n18_), .O(new_n1108_));
  OR       g1092(.a(new_n1108_), .b(new_n1105_), .O(new_n1109_));
  OR       g1093(.a(new_n1109_), .b(new_n1103_), .O(new_n1110_));
  OR       g1094(.a(new_n1110_), .b(new_n1100_), .O(new_n1111_));
  OR       g1095(.a(new_n1111_), .b(new_n1094_), .O(new_n1112_));
  AND      g1096(.a(new_n1112_), .b(new_n22_), .O(new_n1113_));
  AND      g1097(.a(new_n24_), .b(i_2_0_49_0), .O(new_n1114_));
  NOT      g1098(.a(new_n1114_), .O(new_n1115_));
  AND      g1099(.a(new_n159_), .b(i_2_0_109_0), .O(new_n1116_));
  AND      g1100(.a(new_n1116_), .b(new_n1115_), .O(new_n1117_));
  OR       g1101(.a(new_n63_), .b(i_2_0_49_0), .O(new_n1118_));
  NAND     g1102(.a(new_n1118_), .b(new_n176_), .O(new_n1119_));
  OR       g1103(.a(new_n1119_), .b(new_n747_), .O(new_n1120_));
  OR       g1104(.a(new_n1120_), .b(new_n1117_), .O(new_n1121_));
  NAND     g1105(.a(new_n1121_), .b(new_n949_), .O(new_n1122_));
  AND      g1106(.a(new_n1122_), .b(new_n364_), .O(new_n1123_));
  AND      g1107(.a(i_2_0_49_0), .b(i_2_0_16_0), .O(new_n1124_));
  OR       g1108(.a(new_n1009_), .b(new_n444_), .O(new_n1125_));
  AND      g1109(.a(new_n206_), .b(new_n180_), .O(new_n1126_));
  NAND     g1110(.a(new_n992_), .b(new_n135_), .O(new_n1127_));
  OR       g1111(.a(new_n92_), .b(new_n152_), .O(new_n1128_));
  AND      g1112(.a(new_n1128_), .b(new_n1127_), .O(new_n1129_));
  AND      g1113(.a(new_n1129_), .b(new_n1126_), .O(new_n1130_));
  NAND     g1114(.a(new_n1130_), .b(new_n1125_), .O(new_n1131_));
  AND      g1115(.a(new_n1131_), .b(new_n1124_), .O(new_n1132_));
  OR       g1116(.a(new_n1132_), .b(new_n1123_), .O(new_n1133_));
  OR       g1117(.a(new_n1133_), .b(new_n1113_), .O(new_n1134_));
  AND      g1118(.a(new_n1134_), .b(new_n82_), .O(new_n1135_));
  NAND     g1119(.a(new_n754_), .b(new_n426_), .O(new_n1136_));
  AND      g1120(.a(new_n1118_), .b(new_n33_), .O(new_n1137_));
  AND      g1121(.a(new_n1137_), .b(new_n1136_), .O(new_n1138_));
  AND      g1122(.a(new_n34_), .b(i_2_0_109_0), .O(new_n1139_));
  OR       g1123(.a(new_n1139_), .b(new_n1124_), .O(new_n1140_));
  OR       g1124(.a(new_n1140_), .b(new_n1138_), .O(new_n1141_));
  AND      g1125(.a(new_n1141_), .b(i_2_0_66_0), .O(new_n1142_));
  OR       g1126(.a(new_n175_), .b(i_2_0_74_0), .O(new_n1143_));
  NAND     g1127(.a(new_n1143_), .b(new_n97_), .O(new_n1144_));
  AND      g1128(.a(new_n1144_), .b(new_n992_), .O(new_n1145_));
  NAND     g1129(.a(new_n577_), .b(new_n134_), .O(new_n1146_));
  OR       g1130(.a(new_n754_), .b(new_n596_), .O(new_n1147_));
  NAND     g1131(.a(new_n1147_), .b(new_n1146_), .O(new_n1148_));
  AND      g1132(.a(new_n1148_), .b(i_2_0_74_0), .O(new_n1149_));
  OR       g1133(.a(new_n1149_), .b(new_n1145_), .O(new_n1150_));
  AND      g1134(.a(new_n1150_), .b(new_n21_), .O(new_n1151_));
  AND      g1135(.a(new_n83_), .b(new_n65_), .O(new_n1152_));
  OR       g1136(.a(new_n51_), .b(new_n17_), .O(new_n1153_));
  OR       g1137(.a(new_n1153_), .b(new_n710_), .O(new_n1154_));
  OR       g1138(.a(new_n963_), .b(new_n168_), .O(new_n1155_));
  OR       g1139(.a(new_n1155_), .b(new_n248_), .O(new_n1156_));
  NAND     g1140(.a(new_n1156_), .b(new_n1154_), .O(new_n1157_));
  AND      g1141(.a(new_n34_), .b(new_n62_), .O(new_n1158_));
  AND      g1142(.a(new_n283_), .b(new_n64_), .O(new_n1159_));
  OR       g1143(.a(new_n1159_), .b(new_n1158_), .O(new_n1160_));
  OR       g1144(.a(new_n1160_), .b(new_n1157_), .O(new_n1161_));
  OR       g1145(.a(new_n1161_), .b(new_n1152_), .O(new_n1162_));
  AND      g1146(.a(new_n1162_), .b(i_2_0_118_0), .O(new_n1163_));
  OR       g1147(.a(new_n1163_), .b(new_n1151_), .O(new_n1164_));
  OR       g1148(.a(new_n1164_), .b(new_n1142_), .O(new_n1165_));
  AND      g1149(.a(new_n702_), .b(i_2_0_49_0), .O(new_n1166_));
  OR       g1150(.a(new_n1166_), .b(new_n527_), .O(new_n1167_));
  AND      g1151(.a(new_n1167_), .b(new_n1104_), .O(new_n1168_));
  OR       g1152(.a(new_n992_), .b(new_n333_), .O(new_n1169_));
  AND      g1153(.a(new_n1169_), .b(new_n51_), .O(new_n1170_));
  NAND     g1154(.a(new_n477_), .b(i_2_0_109_0), .O(new_n1171_));
  NAND     g1155(.a(new_n1171_), .b(new_n1079_), .O(new_n1172_));
  OR       g1156(.a(new_n1172_), .b(new_n1170_), .O(new_n1173_));
  AND      g1157(.a(new_n1173_), .b(new_n1058_), .O(new_n1174_));
  NOT      g1158(.a(new_n1003_), .O(new_n1175_));
  OR       g1159(.a(new_n661_), .b(new_n164_), .O(new_n1176_));
  NAND     g1160(.a(new_n1176_), .b(new_n1171_), .O(new_n1177_));
  NAND     g1161(.a(new_n1074_), .b(new_n168_), .O(new_n1178_));
  AND      g1162(.a(new_n1178_), .b(new_n152_), .O(new_n1179_));
  OR       g1163(.a(new_n1179_), .b(new_n1177_), .O(new_n1180_));
  AND      g1164(.a(new_n1180_), .b(new_n1175_), .O(new_n1181_));
  OR       g1165(.a(new_n1181_), .b(new_n1174_), .O(new_n1182_));
  OR       g1166(.a(new_n1182_), .b(new_n1168_), .O(new_n1183_));
  OR       g1167(.a(new_n871_), .b(new_n33_), .O(new_n1184_));
  AND      g1168(.a(new_n1184_), .b(i_2_0_66_0), .O(new_n1185_));
  OR       g1169(.a(new_n1185_), .b(new_n323_), .O(new_n1186_));
  AND      g1170(.a(new_n1186_), .b(new_n1039_), .O(new_n1187_));
  OR       g1171(.a(new_n1187_), .b(new_n1183_), .O(new_n1188_));
  OR       g1172(.a(new_n1188_), .b(new_n1165_), .O(new_n1189_));
  AND      g1173(.a(new_n1189_), .b(new_n372_), .O(new_n1190_));
  NAND     g1174(.a(new_n866_), .b(new_n553_), .O(new_n1191_));
  AND      g1175(.a(new_n1191_), .b(new_n923_), .O(new_n1192_));
  AND      g1176(.a(new_n62_), .b(i_2_0_49_0), .O(new_n1193_));
  NAND     g1177(.a(new_n1153_), .b(new_n758_), .O(new_n1194_));
  AND      g1178(.a(new_n1194_), .b(new_n1193_), .O(new_n1195_));
  OR       g1179(.a(new_n1195_), .b(new_n1192_), .O(new_n1196_));
  OR       g1180(.a(new_n1028_), .b(new_n721_), .O(new_n1197_));
  OR       g1181(.a(new_n113_), .b(i_2_0_118_0), .O(new_n1198_));
  OR       g1182(.a(new_n1198_), .b(new_n992_), .O(new_n1199_));
  NAND     g1183(.a(new_n1199_), .b(new_n1197_), .O(new_n1200_));
  OR       g1184(.a(new_n91_), .b(i_2_0_57_0), .O(new_n1201_));
  NAND     g1185(.a(new_n1201_), .b(new_n42_), .O(new_n1202_));
  AND      g1186(.a(new_n1202_), .b(new_n992_), .O(new_n1203_));
  OR       g1187(.a(new_n1203_), .b(new_n1200_), .O(new_n1204_));
  OR       g1188(.a(new_n1204_), .b(new_n1196_), .O(new_n1205_));
  AND      g1189(.a(new_n1205_), .b(new_n779_), .O(new_n1206_));
  AND      g1190(.a(new_n746_), .b(new_n948_), .O(new_n1207_));
  OR       g1191(.a(new_n942_), .b(new_n493_), .O(new_n1208_));
  OR       g1192(.a(new_n1208_), .b(new_n1207_), .O(new_n1209_));
  OR       g1193(.a(new_n1052_), .b(new_n918_), .O(new_n1210_));
  NAND     g1194(.a(new_n1210_), .b(new_n1209_), .O(new_n1211_));
  OR       g1195(.a(new_n1211_), .b(new_n1206_), .O(new_n1212_));
  AND      g1196(.a(new_n1212_), .b(i_2_0_16_0), .O(new_n1213_));
  OR       g1197(.a(new_n1213_), .b(new_n1190_), .O(new_n1214_));
  OR       g1198(.a(new_n1214_), .b(new_n1135_), .O(new_n1215_));
  AND      g1199(.a(new_n1215_), .b(i_2_0_13_0), .O(new_n1216_));
  OR       g1200(.a(new_n138_), .b(new_n41_), .O(new_n1217_));
  NAND     g1201(.a(new_n1217_), .b(new_n766_), .O(new_n1218_));
  AND      g1202(.a(new_n1218_), .b(new_n163_), .O(new_n1219_));
  AND      g1203(.a(new_n98_), .b(new_n33_), .O(new_n1220_));
  AND      g1204(.a(new_n1220_), .b(new_n803_), .O(new_n1221_));
  NAND     g1205(.a(new_n113_), .b(i_2_0_142_0), .O(new_n1222_));
  AND      g1206(.a(new_n1222_), .b(new_n321_), .O(new_n1223_));
  AND      g1207(.a(new_n762_), .b(new_n192_), .O(new_n1224_));
  OR       g1208(.a(new_n1224_), .b(new_n1223_), .O(new_n1225_));
  OR       g1209(.a(new_n1225_), .b(new_n1221_), .O(new_n1226_));
  OR       g1210(.a(new_n1226_), .b(new_n1219_), .O(new_n1227_));
  AND      g1211(.a(new_n1227_), .b(i_2_0_49_0), .O(new_n1228_));
  OR       g1212(.a(new_n1139_), .b(new_n503_), .O(new_n1229_));
  AND      g1213(.a(new_n1229_), .b(new_n585_), .O(new_n1230_));
  OR       g1214(.a(new_n1106_), .b(new_n22_), .O(new_n1231_));
  AND      g1215(.a(new_n678_), .b(new_n63_), .O(new_n1232_));
  AND      g1216(.a(new_n1232_), .b(new_n1231_), .O(new_n1233_));
  OR       g1217(.a(new_n1233_), .b(new_n1230_), .O(new_n1234_));
  OR       g1218(.a(new_n1234_), .b(new_n1228_), .O(new_n1235_));
  AND      g1219(.a(new_n1124_), .b(new_n21_), .O(new_n1236_));
  OR       g1220(.a(new_n1236_), .b(new_n264_), .O(new_n1237_));
  OR       g1221(.a(i_2_0_49_0), .b(i_2_0_16_0), .O(new_n1238_));
  AND      g1222(.a(new_n1238_), .b(i_2_0_66_0), .O(new_n1239_));
  AND      g1223(.a(new_n1239_), .b(new_n1237_), .O(new_n1240_));
  AND      g1224(.a(new_n762_), .b(new_n25_), .O(new_n1241_));
  AND      g1225(.a(new_n503_), .b(new_n21_), .O(new_n1242_));
  OR       g1226(.a(new_n1059_), .b(new_n82_), .O(new_n1243_));
  AND      g1227(.a(new_n1243_), .b(new_n1242_), .O(new_n1244_));
  OR       g1228(.a(new_n1244_), .b(new_n1241_), .O(new_n1245_));
  OR       g1229(.a(new_n1245_), .b(new_n1240_), .O(new_n1246_));
  AND      g1230(.a(new_n1246_), .b(new_n152_), .O(new_n1247_));
  OR       g1231(.a(new_n1247_), .b(new_n1235_), .O(new_n1248_));
  AND      g1232(.a(new_n1248_), .b(new_n419_), .O(new_n1249_));
  NAND     g1233(.a(new_n1058_), .b(new_n265_), .O(new_n1250_));
  NAND     g1234(.a(new_n34_), .b(new_n29_), .O(new_n1251_));
  OR       g1235(.a(new_n1251_), .b(new_n493_), .O(new_n1252_));
  NAND     g1236(.a(new_n1252_), .b(new_n1250_), .O(new_n1253_));
  AND      g1237(.a(new_n1253_), .b(new_n63_), .O(new_n1254_));
  OR       g1238(.a(new_n1114_), .b(new_n34_), .O(new_n1255_));
  AND      g1239(.a(new_n372_), .b(new_n69_), .O(new_n1256_));
  AND      g1240(.a(new_n1256_), .b(new_n1255_), .O(new_n1257_));
  AND      g1241(.a(new_n1106_), .b(new_n638_), .O(new_n1258_));
  NAND     g1242(.a(new_n778_), .b(i_2_0_142_0), .O(new_n1259_));
  AND      g1243(.a(new_n1259_), .b(new_n1058_), .O(new_n1260_));
  OR       g1244(.a(new_n1260_), .b(new_n372_), .O(new_n1261_));
  OR       g1245(.a(new_n1261_), .b(new_n1258_), .O(new_n1262_));
  AND      g1246(.a(new_n1262_), .b(new_n22_), .O(new_n1263_));
  OR       g1247(.a(new_n1263_), .b(new_n1257_), .O(new_n1264_));
  OR       g1248(.a(new_n1264_), .b(new_n1254_), .O(new_n1265_));
  AND      g1249(.a(new_n1265_), .b(i_2_0_66_0), .O(new_n1266_));
  NAND     g1250(.a(new_n785_), .b(new_n383_), .O(new_n1267_));
  AND      g1251(.a(new_n1124_), .b(new_n321_), .O(new_n1268_));
  AND      g1252(.a(new_n1268_), .b(new_n1267_), .O(new_n1269_));
  NAND     g1253(.a(new_n1236_), .b(new_n372_), .O(new_n1270_));
  OR       g1254(.a(new_n383_), .b(new_n753_), .O(new_n1271_));
  AND      g1255(.a(new_n1271_), .b(new_n29_), .O(new_n1272_));
  OR       g1256(.a(new_n1077_), .b(new_n367_), .O(new_n1273_));
  OR       g1257(.a(new_n1273_), .b(new_n1272_), .O(new_n1274_));
  NAND     g1258(.a(new_n1274_), .b(new_n1270_), .O(new_n1275_));
  OR       g1259(.a(new_n1275_), .b(new_n1269_), .O(new_n1276_));
  OR       g1260(.a(new_n1276_), .b(new_n1266_), .O(new_n1277_));
  OR       g1261(.a(new_n1238_), .b(new_n401_), .O(new_n1278_));
  AND      g1262(.a(new_n1278_), .b(new_n82_), .O(new_n1279_));
  OR       g1263(.a(new_n1279_), .b(new_n1236_), .O(new_n1280_));
  AND      g1264(.a(new_n1280_), .b(new_n638_), .O(new_n1281_));
  OR       g1265(.a(new_n28_), .b(new_n77_), .O(new_n1282_));
  OR       g1266(.a(new_n1282_), .b(new_n1074_), .O(new_n1283_));
  AND      g1267(.a(new_n391_), .b(new_n77_), .O(new_n1284_));
  OR       g1268(.a(new_n1284_), .b(new_n44_), .O(new_n1285_));
  NAND     g1269(.a(new_n1285_), .b(new_n1283_), .O(new_n1286_));
  OR       g1270(.a(new_n1286_), .b(new_n1281_), .O(new_n1287_));
  AND      g1271(.a(new_n564_), .b(new_n110_), .O(new_n1288_));
  NAND     g1272(.a(new_n1288_), .b(new_n384_), .O(new_n1289_));
  AND      g1273(.a(new_n1289_), .b(new_n1124_), .O(new_n1290_));
  AND      g1274(.a(new_n790_), .b(new_n135_), .O(new_n1291_));
  OR       g1275(.a(new_n137_), .b(new_n753_), .O(new_n1292_));
  NAND     g1276(.a(new_n1292_), .b(new_n785_), .O(new_n1293_));
  OR       g1277(.a(new_n1293_), .b(new_n1291_), .O(new_n1294_));
  OR       g1278(.a(new_n1236_), .b(new_n19_), .O(new_n1295_));
  AND      g1279(.a(new_n1295_), .b(new_n662_), .O(new_n1296_));
  AND      g1280(.a(new_n1296_), .b(new_n1294_), .O(new_n1297_));
  OR       g1281(.a(new_n1297_), .b(new_n1290_), .O(new_n1298_));
  OR       g1282(.a(new_n1298_), .b(new_n1287_), .O(new_n1299_));
  AND      g1283(.a(new_n1299_), .b(new_n63_), .O(new_n1300_));
  NAND     g1284(.a(new_n835_), .b(new_n45_), .O(new_n1301_));
  AND      g1285(.a(new_n1301_), .b(new_n520_), .O(new_n1302_));
  OR       g1286(.a(new_n44_), .b(new_n97_), .O(new_n1303_));
  OR       g1287(.a(new_n485_), .b(new_n54_), .O(new_n1304_));
  NAND     g1288(.a(new_n1304_), .b(new_n1303_), .O(new_n1305_));
  OR       g1289(.a(new_n1305_), .b(new_n1302_), .O(new_n1306_));
  AND      g1290(.a(new_n1306_), .b(i_2_0_49_0), .O(new_n1307_));
  OR       g1291(.a(new_n778_), .b(new_n24_), .O(new_n1308_));
  NAND     g1292(.a(new_n1308_), .b(new_n105_), .O(new_n1309_));
  AND      g1293(.a(new_n1309_), .b(new_n1175_), .O(new_n1310_));
  AND      g1294(.a(new_n1101_), .b(new_n98_), .O(new_n1311_));
  AND      g1295(.a(new_n1311_), .b(new_n265_), .O(new_n1312_));
  OR       g1296(.a(new_n1282_), .b(new_n683_), .O(new_n1313_));
  OR       g1297(.a(new_n107_), .b(i_2_0_139_0), .O(new_n1314_));
  OR       g1298(.a(new_n1314_), .b(new_n1251_), .O(new_n1315_));
  NAND     g1299(.a(new_n1315_), .b(new_n1313_), .O(new_n1316_));
  OR       g1300(.a(new_n1316_), .b(new_n1312_), .O(new_n1317_));
  OR       g1301(.a(new_n1317_), .b(new_n1310_), .O(new_n1318_));
  OR       g1302(.a(new_n1318_), .b(new_n1307_), .O(new_n1319_));
  AND      g1303(.a(new_n1319_), .b(new_n924_), .O(new_n1320_));
  OR       g1304(.a(new_n1320_), .b(new_n1300_), .O(new_n1321_));
  OR       g1305(.a(new_n1321_), .b(new_n1277_), .O(new_n1322_));
  NAND     g1306(.a(new_n28_), .b(new_n92_), .O(new_n1323_));
  AND      g1307(.a(new_n1323_), .b(new_n1058_), .O(new_n1324_));
  OR       g1308(.a(new_n54_), .b(i_2_0_118_0), .O(new_n1325_));
  NAND     g1309(.a(new_n1325_), .b(new_n188_), .O(new_n1326_));
  OR       g1310(.a(new_n1326_), .b(new_n1324_), .O(new_n1327_));
  AND      g1311(.a(new_n1327_), .b(new_n22_), .O(new_n1328_));
  NAND     g1312(.a(new_n1271_), .b(new_n54_), .O(new_n1329_));
  AND      g1313(.a(new_n1329_), .b(new_n64_), .O(new_n1330_));
  OR       g1314(.a(new_n188_), .b(new_n24_), .O(new_n1331_));
  OR       g1315(.a(new_n383_), .b(new_n121_), .O(new_n1332_));
  NAND     g1316(.a(new_n1332_), .b(new_n1331_), .O(new_n1333_));
  AND      g1317(.a(new_n803_), .b(new_n41_), .O(new_n1334_));
  AND      g1318(.a(new_n1334_), .b(new_n1333_), .O(new_n1335_));
  OR       g1319(.a(new_n1335_), .b(new_n1330_), .O(new_n1336_));
  OR       g1320(.a(new_n1336_), .b(new_n1328_), .O(new_n1337_));
  AND      g1321(.a(new_n1337_), .b(new_n152_), .O(new_n1338_));
  AND      g1322(.a(new_n803_), .b(new_n303_), .O(new_n1339_));
  AND      g1323(.a(new_n82_), .b(i_2_0_49_0), .O(new_n1340_));
  NAND     g1324(.a(new_n1003_), .b(new_n41_), .O(new_n1341_));
  AND      g1325(.a(new_n1341_), .b(new_n1340_), .O(new_n1342_));
  OR       g1326(.a(new_n1342_), .b(new_n1339_), .O(new_n1343_));
  AND      g1327(.a(new_n1343_), .b(new_n1106_), .O(new_n1344_));
  NOT      g1328(.a(new_n803_), .O(new_n1345_));
  NAND     g1329(.a(new_n1002_), .b(new_n1345_), .O(new_n1346_));
  AND      g1330(.a(new_n1346_), .b(new_n1078_), .O(new_n1347_));
  NAND     g1331(.a(i_2_0_143_0), .b(i_2_0_118_0), .O(new_n1348_));
  NAND     g1332(.a(new_n1348_), .b(new_n963_), .O(new_n1349_));
  AND      g1333(.a(new_n1349_), .b(new_n177_), .O(new_n1350_));
  AND      g1334(.a(new_n1350_), .b(new_n1139_), .O(new_n1351_));
  OR       g1335(.a(new_n1351_), .b(new_n1347_), .O(new_n1352_));
  OR       g1336(.a(new_n1352_), .b(new_n1344_), .O(new_n1353_));
  OR       g1337(.a(new_n107_), .b(i_2_0_49_0), .O(new_n1354_));
  AND      g1338(.a(new_n1354_), .b(new_n1115_), .O(new_n1355_));
  OR       g1339(.a(new_n1355_), .b(new_n1011_), .O(new_n1356_));
  NAND     g1340(.a(new_n1356_), .b(new_n43_), .O(new_n1357_));
  AND      g1341(.a(new_n1357_), .b(new_n756_), .O(new_n1358_));
  OR       g1342(.a(new_n1358_), .b(new_n1353_), .O(new_n1359_));
  OR       g1343(.a(new_n1359_), .b(new_n1338_), .O(new_n1360_));
  AND      g1344(.a(new_n1360_), .b(new_n62_), .O(new_n1361_));
  OR       g1345(.a(new_n1361_), .b(new_n1322_), .O(new_n1362_));
  OR       g1346(.a(new_n1362_), .b(new_n1249_), .O(new_n1363_));
  AND      g1347(.a(new_n1363_), .b(new_n294_), .O(new_n1364_));
  OR       g1348(.a(new_n1364_), .b(new_n1216_), .O(new_n1365_));
  OR       g1349(.a(new_n1365_), .b(new_n1085_), .O(new_n1366_));
  OR       g1350(.a(new_n1366_), .b(new_n903_), .O(o_2_0_0_0));
endmodule


