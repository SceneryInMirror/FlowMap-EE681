// Benchmark "kernel_2_2" written by ABC on Wed May  4 16:42:25 2022

module kernel_2_2 ( 
    i_2_2_43_0, i_2_2_58_0, i_2_2_60_0, i_2_2_63_0, i_2_2_82_0, i_2_2_91_0,
    i_2_2_107_0, i_2_2_108_0, i_2_2_113_0, i_2_2_116_0, i_2_2_129_0,
    i_2_2_134_0, i_2_2_137_0, i_2_2_139_0, i_2_2_147_0,
    o_2_2_0_0  );
  input  i_2_2_43_0, i_2_2_58_0, i_2_2_60_0, i_2_2_63_0, i_2_2_82_0,
    i_2_2_91_0, i_2_2_107_0, i_2_2_108_0, i_2_2_113_0, i_2_2_116_0,
    i_2_2_129_0, i_2_2_134_0, i_2_2_137_0, i_2_2_139_0, i_2_2_147_0;
  output o_2_2_0_0;
  wire new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_;
  NOT      g000(.a(i_2_2_113_0), .O(new_n17_));
  NOT      g001(.a(i_2_2_108_0), .O(new_n18_));
  NOT      g002(.a(i_2_2_147_0), .O(new_n19_));
  NOT      g003(.a(i_2_2_60_0), .O(new_n20_));
  NOT      g004(.a(i_2_2_107_0), .O(new_n21_));
  OR       g005(.a(i_2_2_137_0), .b(i_2_2_134_0), .O(new_n22_));
  AND      g006(.a(i_2_2_139_0), .b(i_2_2_129_0), .O(new_n23_));
  NOT      g007(.a(new_n23_), .O(new_n24_));
  OR       g008(.a(new_n24_), .b(new_n22_), .O(new_n25_));
  OR       g009(.a(new_n25_), .b(new_n21_), .O(new_n26_));
  AND      g010(.a(i_2_2_137_0), .b(i_2_2_134_0), .O(new_n27_));
  AND      g011(.a(new_n27_), .b(new_n21_), .O(new_n28_));
  NOT      g012(.a(new_n28_), .O(new_n29_));
  NAND     g013(.a(new_n29_), .b(new_n26_), .O(new_n30_));
  AND      g014(.a(new_n30_), .b(i_2_2_91_0), .O(new_n31_));
  AND      g015(.a(new_n23_), .b(i_2_2_137_0), .O(new_n32_));
  AND      g016(.a(new_n32_), .b(i_2_2_134_0), .O(new_n33_));
  OR       g017(.a(new_n33_), .b(new_n31_), .O(new_n34_));
  AND      g018(.a(new_n34_), .b(i_2_2_58_0), .O(new_n35_));
  AND      g019(.a(new_n28_), .b(i_2_2_129_0), .O(new_n36_));
  OR       g020(.a(new_n36_), .b(new_n35_), .O(new_n37_));
  AND      g021(.a(new_n37_), .b(new_n20_), .O(new_n38_));
  NOT      g022(.a(i_2_2_82_0), .O(new_n39_));
  NOT      g023(.a(i_2_2_91_0), .O(new_n40_));
  NOT      g024(.a(i_2_2_137_0), .O(new_n41_));
  OR       g025(.a(i_2_2_139_0), .b(i_2_2_129_0), .O(new_n42_));
  NAND     g026(.a(new_n42_), .b(new_n41_), .O(new_n43_));
  AND      g027(.a(i_2_2_139_0), .b(i_2_2_134_0), .O(new_n44_));
  OR       g028(.a(i_2_2_107_0), .b(i_2_2_58_0), .O(new_n45_));
  OR       g029(.a(new_n45_), .b(new_n44_), .O(new_n46_));
  OR       g030(.a(new_n46_), .b(new_n43_), .O(new_n47_));
  NOT      g031(.a(i_2_2_129_0), .O(new_n48_));
  OR       g032(.a(i_2_2_139_0), .b(new_n48_), .O(new_n49_));
  AND      g033(.a(i_2_2_134_0), .b(i_2_2_58_0), .O(new_n50_));
  NAND     g034(.a(new_n50_), .b(new_n49_), .O(new_n51_));
  AND      g035(.a(new_n51_), .b(new_n47_), .O(new_n52_));
  OR       g036(.a(new_n52_), .b(new_n40_), .O(new_n53_));
  NOT      g037(.a(i_2_2_58_0), .O(new_n54_));
  AND      g038(.a(i_2_2_129_0), .b(new_n21_), .O(new_n55_));
  NAND     g039(.a(new_n55_), .b(i_2_2_134_0), .O(new_n56_));
  OR       g040(.a(new_n56_), .b(new_n54_), .O(new_n57_));
  NAND     g041(.a(new_n57_), .b(new_n53_), .O(new_n58_));
  AND      g042(.a(new_n58_), .b(new_n20_), .O(new_n59_));
  NOT      g043(.a(i_2_2_134_0), .O(new_n60_));
  OR       g044(.a(i_2_2_139_0), .b(new_n60_), .O(new_n61_));
  NOT      g045(.a(i_2_2_139_0), .O(new_n62_));
  OR       g046(.a(new_n62_), .b(i_2_2_107_0), .O(new_n63_));
  OR       g047(.a(new_n63_), .b(i_2_2_91_0), .O(new_n64_));
  NAND     g048(.a(new_n64_), .b(new_n61_), .O(new_n65_));
  AND      g049(.a(new_n65_), .b(i_2_2_129_0), .O(new_n66_));
  OR       g050(.a(i_2_2_129_0), .b(i_2_2_91_0), .O(new_n67_));
  NAND     g051(.a(new_n67_), .b(new_n63_), .O(new_n68_));
  AND      g052(.a(new_n68_), .b(i_2_2_134_0), .O(new_n69_));
  OR       g053(.a(new_n69_), .b(new_n66_), .O(new_n70_));
  AND      g054(.a(new_n70_), .b(i_2_2_137_0), .O(new_n71_));
  AND      g055(.a(i_2_2_91_0), .b(i_2_2_58_0), .O(new_n72_));
  NOT      g056(.a(new_n72_), .O(new_n73_));
  OR       g057(.a(new_n73_), .b(new_n25_), .O(new_n74_));
  OR       g058(.a(new_n41_), .b(i_2_2_129_0), .O(new_n75_));
  OR       g059(.a(new_n75_), .b(new_n73_), .O(new_n76_));
  NAND     g060(.a(new_n44_), .b(i_2_2_129_0), .O(new_n77_));
  OR       g061(.a(new_n77_), .b(new_n45_), .O(new_n78_));
  AND      g062(.a(new_n78_), .b(new_n76_), .O(new_n79_));
  OR       g063(.a(new_n79_), .b(new_n20_), .O(new_n80_));
  NAND     g064(.a(new_n80_), .b(new_n74_), .O(new_n81_));
  OR       g065(.a(new_n81_), .b(new_n71_), .O(new_n82_));
  OR       g066(.a(new_n82_), .b(new_n59_), .O(new_n83_));
  AND      g067(.a(new_n83_), .b(new_n39_), .O(new_n84_));
  AND      g068(.a(i_2_2_82_0), .b(i_2_2_60_0), .O(new_n85_));
  AND      g069(.a(new_n85_), .b(new_n72_), .O(new_n86_));
  AND      g070(.a(new_n86_), .b(new_n32_), .O(new_n87_));
  OR       g071(.a(new_n87_), .b(new_n84_), .O(new_n88_));
  OR       g072(.a(new_n88_), .b(new_n38_), .O(new_n89_));
  AND      g073(.a(new_n89_), .b(i_2_2_63_0), .O(new_n90_));
  AND      g074(.a(i_2_2_129_0), .b(i_2_2_91_0), .O(new_n91_));
  AND      g075(.a(new_n91_), .b(new_n28_), .O(new_n92_));
  NOT      g076(.a(new_n27_), .O(new_n93_));
  OR       g077(.a(i_2_2_107_0), .b(new_n40_), .O(new_n94_));
  OR       g078(.a(new_n94_), .b(new_n62_), .O(new_n95_));
  OR       g079(.a(new_n95_), .b(new_n48_), .O(new_n96_));
  NAND     g080(.a(new_n96_), .b(new_n93_), .O(new_n97_));
  OR       g081(.a(i_2_2_82_0), .b(i_2_2_60_0), .O(new_n98_));
  NOT      g082(.a(new_n98_), .O(new_n99_));
  AND      g083(.a(new_n99_), .b(new_n22_), .O(new_n100_));
  AND      g084(.a(new_n100_), .b(new_n97_), .O(new_n101_));
  OR       g085(.a(new_n101_), .b(new_n92_), .O(new_n102_));
  NOT      g086(.a(new_n85_), .O(new_n103_));
  AND      g087(.a(new_n103_), .b(i_2_2_58_0), .O(new_n104_));
  AND      g088(.a(new_n104_), .b(new_n102_), .O(new_n105_));
  OR       g089(.a(new_n105_), .b(new_n90_), .O(new_n106_));
  AND      g090(.a(new_n106_), .b(i_2_2_116_0), .O(new_n107_));
  NOT      g091(.a(i_2_2_116_0), .O(new_n108_));
  AND      g092(.a(new_n108_), .b(i_2_2_91_0), .O(new_n109_));
  NAND     g093(.a(new_n109_), .b(i_2_2_137_0), .O(new_n110_));
  XOR      g094(.a(i_2_2_137_0), .b(new_n60_), .O(new_n111_));
  AND      g095(.a(i_2_2_129_0), .b(i_2_2_58_0), .O(new_n112_));
  NAND     g096(.a(new_n112_), .b(new_n111_), .O(new_n113_));
  AND      g097(.a(new_n113_), .b(new_n110_), .O(new_n114_));
  NOT      g098(.a(i_2_2_63_0), .O(new_n115_));
  AND      g099(.a(new_n63_), .b(new_n60_), .O(new_n116_));
  OR       g100(.a(new_n116_), .b(new_n115_), .O(new_n117_));
  OR       g101(.a(new_n117_), .b(new_n114_), .O(new_n118_));
  AND      g102(.a(new_n27_), .b(i_2_2_139_0), .O(new_n119_));
  NAND     g103(.a(new_n119_), .b(new_n109_), .O(new_n120_));
  NAND     g104(.a(new_n120_), .b(new_n118_), .O(new_n121_));
  AND      g105(.a(new_n121_), .b(new_n39_), .O(new_n122_));
  NOT      g106(.a(new_n95_), .O(new_n123_));
  OR       g107(.a(i_2_2_129_0), .b(i_2_2_116_0), .O(new_n124_));
  NOT      g108(.a(new_n124_), .O(new_n125_));
  AND      g109(.a(new_n125_), .b(new_n27_), .O(new_n126_));
  AND      g110(.a(new_n126_), .b(new_n123_), .O(new_n127_));
  OR       g111(.a(new_n127_), .b(new_n122_), .O(new_n128_));
  AND      g112(.a(new_n128_), .b(new_n20_), .O(new_n129_));
  OR       g113(.a(new_n129_), .b(new_n107_), .O(new_n130_));
  AND      g114(.a(new_n130_), .b(new_n19_), .O(new_n131_));
  AND      g115(.a(i_2_2_116_0), .b(new_n21_), .O(new_n132_));
  AND      g116(.a(new_n132_), .b(i_2_2_58_0), .O(new_n133_));
  AND      g117(.a(i_2_2_129_0), .b(i_2_2_63_0), .O(new_n134_));
  AND      g118(.a(new_n134_), .b(new_n109_), .O(new_n135_));
  OR       g119(.a(new_n135_), .b(new_n133_), .O(new_n136_));
  AND      g120(.a(new_n136_), .b(i_2_2_139_0), .O(new_n137_));
  AND      g121(.a(new_n62_), .b(i_2_2_91_0), .O(new_n138_));
  AND      g122(.a(new_n138_), .b(new_n134_), .O(new_n139_));
  OR       g123(.a(new_n91_), .b(i_2_2_63_0), .O(new_n140_));
  AND      g124(.a(new_n21_), .b(i_2_2_58_0), .O(new_n141_));
  AND      g125(.a(new_n141_), .b(new_n140_), .O(new_n142_));
  OR       g126(.a(new_n142_), .b(new_n139_), .O(new_n143_));
  AND      g127(.a(new_n143_), .b(i_2_2_116_0), .O(new_n144_));
  OR       g128(.a(new_n144_), .b(new_n137_), .O(new_n145_));
  AND      g129(.a(new_n145_), .b(new_n20_), .O(new_n146_));
  AND      g130(.a(i_2_2_116_0), .b(i_2_2_91_0), .O(new_n147_));
  AND      g131(.a(i_2_2_139_0), .b(i_2_2_63_0), .O(new_n148_));
  AND      g132(.a(new_n148_), .b(new_n147_), .O(new_n149_));
  AND      g133(.a(new_n149_), .b(new_n112_), .O(new_n150_));
  OR       g134(.a(new_n150_), .b(new_n146_), .O(new_n151_));
  AND      g135(.a(i_2_2_134_0), .b(new_n39_), .O(new_n152_));
  AND      g136(.a(new_n152_), .b(i_2_2_137_0), .O(new_n153_));
  AND      g137(.a(new_n153_), .b(new_n151_), .O(new_n154_));
  OR       g138(.a(new_n154_), .b(new_n131_), .O(new_n155_));
  AND      g139(.a(new_n155_), .b(new_n18_), .O(new_n156_));
  NOT      g140(.a(i_2_2_43_0), .O(new_n157_));
  NAND     g141(.a(i_2_2_116_0), .b(i_2_2_91_0), .O(new_n158_));
  OR       g142(.a(i_2_2_107_0), .b(i_2_2_82_0), .O(new_n159_));
  NAND     g143(.a(new_n159_), .b(new_n158_), .O(new_n160_));
  AND      g144(.a(new_n160_), .b(new_n42_), .O(new_n161_));
  OR       g145(.a(new_n161_), .b(new_n132_), .O(new_n162_));
  AND      g146(.a(new_n162_), .b(i_2_2_63_0), .O(new_n163_));
  OR       g147(.a(new_n95_), .b(new_n108_), .O(new_n164_));
  AND      g148(.a(new_n94_), .b(new_n108_), .O(new_n165_));
  OR       g149(.a(new_n165_), .b(i_2_2_82_0), .O(new_n166_));
  OR       g150(.a(new_n166_), .b(new_n125_), .O(new_n167_));
  NAND     g151(.a(new_n167_), .b(new_n164_), .O(new_n168_));
  OR       g152(.a(new_n168_), .b(new_n163_), .O(new_n169_));
  AND      g153(.a(new_n169_), .b(i_2_2_58_0), .O(new_n170_));
  OR       g154(.a(new_n21_), .b(i_2_2_63_0), .O(new_n171_));
  AND      g155(.a(new_n171_), .b(i_2_2_116_0), .O(new_n172_));
  AND      g156(.a(new_n21_), .b(i_2_2_63_0), .O(new_n173_));
  NAND     g157(.a(new_n173_), .b(i_2_2_139_0), .O(new_n174_));
  NAND     g158(.a(new_n174_), .b(i_2_2_82_0), .O(new_n175_));
  OR       g159(.a(new_n175_), .b(new_n172_), .O(new_n176_));
  OR       g160(.a(i_2_2_129_0), .b(new_n40_), .O(new_n177_));
  OR       g161(.a(new_n177_), .b(i_2_2_139_0), .O(new_n178_));
  AND      g162(.a(new_n178_), .b(i_2_2_116_0), .O(new_n179_));
  AND      g163(.a(new_n91_), .b(i_2_2_139_0), .O(new_n180_));
  AND      g164(.a(new_n180_), .b(new_n171_), .O(new_n181_));
  OR       g165(.a(new_n181_), .b(new_n179_), .O(new_n182_));
  OR       g166(.a(new_n182_), .b(new_n176_), .O(new_n183_));
  AND      g167(.a(new_n183_), .b(new_n19_), .O(new_n184_));
  OR       g168(.a(new_n184_), .b(new_n170_), .O(new_n185_));
  NAND     g169(.a(new_n95_), .b(new_n108_), .O(new_n186_));
  AND      g170(.a(new_n186_), .b(i_2_2_63_0), .O(new_n187_));
  OR       g171(.a(new_n134_), .b(i_2_2_116_0), .O(new_n188_));
  AND      g172(.a(i_2_2_139_0), .b(new_n21_), .O(new_n189_));
  OR       g173(.a(new_n138_), .b(new_n189_), .O(new_n190_));
  AND      g174(.a(new_n190_), .b(new_n188_), .O(new_n191_));
  OR       g175(.a(new_n191_), .b(new_n187_), .O(new_n192_));
  AND      g176(.a(new_n192_), .b(new_n39_), .O(new_n193_));
  OR       g177(.a(new_n94_), .b(i_2_2_139_0), .O(new_n194_));
  NAND     g178(.a(new_n194_), .b(new_n174_), .O(new_n195_));
  AND      g179(.a(new_n195_), .b(new_n179_), .O(new_n196_));
  OR       g180(.a(new_n196_), .b(i_2_2_58_0), .O(new_n197_));
  OR       g181(.a(new_n197_), .b(new_n193_), .O(new_n198_));
  AND      g182(.a(new_n198_), .b(new_n185_), .O(new_n199_));
  OR       g183(.a(new_n42_), .b(i_2_2_91_0), .O(new_n200_));
  AND      g184(.a(new_n200_), .b(i_2_2_63_0), .O(new_n201_));
  OR       g185(.a(new_n201_), .b(new_n180_), .O(new_n202_));
  AND      g186(.a(i_2_2_116_0), .b(new_n39_), .O(new_n203_));
  NAND     g187(.a(new_n94_), .b(new_n48_), .O(new_n204_));
  AND      g188(.a(new_n204_), .b(new_n203_), .O(new_n205_));
  AND      g189(.a(new_n205_), .b(new_n202_), .O(new_n206_));
  OR       g190(.a(new_n206_), .b(new_n199_), .O(new_n207_));
  AND      g191(.a(new_n207_), .b(new_n20_), .O(new_n208_));
  AND      g192(.a(new_n39_), .b(i_2_2_63_0), .O(new_n209_));
  OR       g193(.a(new_n209_), .b(new_n23_), .O(new_n210_));
  AND      g194(.a(new_n210_), .b(i_2_2_91_0), .O(new_n211_));
  OR       g195(.a(i_2_2_139_0), .b(new_n39_), .O(new_n212_));
  OR       g196(.a(new_n212_), .b(new_n134_), .O(new_n213_));
  AND      g197(.a(new_n213_), .b(i_2_2_58_0), .O(new_n214_));
  AND      g198(.a(new_n124_), .b(new_n49_), .O(new_n215_));
  OR       g199(.a(new_n209_), .b(new_n48_), .O(new_n216_));
  AND      g200(.a(new_n216_), .b(new_n215_), .O(new_n217_));
  OR       g201(.a(new_n217_), .b(new_n214_), .O(new_n218_));
  OR       g202(.a(new_n218_), .b(new_n211_), .O(new_n219_));
  AND      g203(.a(new_n219_), .b(new_n19_), .O(new_n220_));
  AND      g204(.a(new_n39_), .b(i_2_2_58_0), .O(new_n221_));
  NAND     g205(.a(new_n42_), .b(new_n115_), .O(new_n222_));
  OR       g206(.a(new_n222_), .b(new_n23_), .O(new_n223_));
  AND      g207(.a(new_n223_), .b(new_n221_), .O(new_n224_));
  OR       g208(.a(new_n224_), .b(new_n220_), .O(new_n225_));
  AND      g209(.a(new_n225_), .b(i_2_2_137_0), .O(new_n226_));
  AND      g210(.a(new_n19_), .b(i_2_2_58_0), .O(new_n227_));
  AND      g211(.a(new_n42_), .b(i_2_2_116_0), .O(new_n228_));
  AND      g212(.a(new_n228_), .b(new_n227_), .O(new_n229_));
  AND      g213(.a(new_n229_), .b(new_n140_), .O(new_n230_));
  OR       g214(.a(new_n230_), .b(new_n226_), .O(new_n231_));
  AND      g215(.a(new_n231_), .b(new_n21_), .O(new_n232_));
  AND      g216(.a(i_2_2_137_0), .b(i_2_2_63_0), .O(new_n233_));
  OR       g217(.a(new_n19_), .b(i_2_2_63_0), .O(new_n234_));
  AND      g218(.a(new_n234_), .b(new_n221_), .O(new_n235_));
  OR       g219(.a(new_n235_), .b(new_n233_), .O(new_n236_));
  AND      g220(.a(new_n236_), .b(i_2_2_116_0), .O(new_n237_));
  AND      g221(.a(new_n19_), .b(i_2_2_137_0), .O(new_n238_));
  AND      g222(.a(new_n238_), .b(new_n221_), .O(new_n239_));
  OR       g223(.a(new_n239_), .b(new_n237_), .O(new_n240_));
  AND      g224(.a(new_n240_), .b(i_2_2_139_0), .O(new_n241_));
  OR       g225(.a(new_n203_), .b(new_n148_), .O(new_n242_));
  OR       g226(.a(i_2_2_116_0), .b(new_n39_), .O(new_n243_));
  AND      g227(.a(new_n243_), .b(new_n227_), .O(new_n244_));
  AND      g228(.a(new_n244_), .b(new_n242_), .O(new_n245_));
  OR       g229(.a(i_2_2_82_0), .b(new_n54_), .O(new_n246_));
  OR       g230(.a(i_2_2_147_0), .b(i_2_2_116_0), .O(new_n247_));
  OR       g231(.a(new_n247_), .b(new_n115_), .O(new_n248_));
  NAND     g232(.a(new_n248_), .b(new_n246_), .O(new_n249_));
  AND      g233(.a(new_n62_), .b(i_2_2_137_0), .O(new_n250_));
  AND      g234(.a(new_n250_), .b(new_n249_), .O(new_n251_));
  OR       g235(.a(new_n251_), .b(new_n245_), .O(new_n252_));
  AND      g236(.a(new_n252_), .b(i_2_2_91_0), .O(new_n253_));
  OR       g237(.a(new_n253_), .b(new_n241_), .O(new_n254_));
  AND      g238(.a(new_n254_), .b(i_2_2_129_0), .O(new_n255_));
  OR       g239(.a(i_2_2_147_0), .b(i_2_2_82_0), .O(new_n256_));
  NOT      g240(.a(new_n256_), .O(new_n257_));
  AND      g241(.a(i_2_2_137_0), .b(i_2_2_116_0), .O(new_n258_));
  AND      g242(.a(new_n258_), .b(new_n257_), .O(new_n259_));
  AND      g243(.a(i_2_2_139_0), .b(i_2_2_137_0), .O(new_n260_));
  OR       g244(.a(new_n260_), .b(new_n147_), .O(new_n261_));
  AND      g245(.a(new_n261_), .b(new_n209_), .O(new_n262_));
  OR       g246(.a(new_n258_), .b(new_n209_), .O(new_n263_));
  OR       g247(.a(i_2_2_137_0), .b(i_2_2_116_0), .O(new_n264_));
  AND      g248(.a(new_n264_), .b(new_n19_), .O(new_n265_));
  AND      g249(.a(new_n265_), .b(new_n263_), .O(new_n266_));
  OR       g250(.a(new_n266_), .b(new_n262_), .O(new_n267_));
  AND      g251(.a(new_n267_), .b(i_2_2_58_0), .O(new_n268_));
  OR       g252(.a(new_n268_), .b(new_n259_), .O(new_n269_));
  OR       g253(.a(new_n269_), .b(new_n255_), .O(new_n270_));
  OR       g254(.a(new_n270_), .b(new_n232_), .O(new_n271_));
  OR       g255(.a(new_n271_), .b(new_n208_), .O(new_n272_));
  AND      g256(.a(new_n272_), .b(i_2_2_134_0), .O(new_n273_));
  AND      g257(.a(new_n67_), .b(i_2_2_63_0), .O(new_n274_));
  OR       g258(.a(new_n274_), .b(i_2_2_129_0), .O(new_n275_));
  AND      g259(.a(new_n238_), .b(new_n133_), .O(new_n276_));
  AND      g260(.a(new_n276_), .b(new_n275_), .O(new_n277_));
  OR       g261(.a(new_n277_), .b(new_n273_), .O(new_n278_));
  NAND     g262(.a(i_2_2_147_0), .b(i_2_2_107_0), .O(new_n279_));
  AND      g263(.a(new_n42_), .b(i_2_2_91_0), .O(new_n280_));
  OR       g264(.a(new_n280_), .b(new_n279_), .O(new_n281_));
  AND      g265(.a(new_n281_), .b(i_2_2_116_0), .O(new_n282_));
  OR       g266(.a(new_n282_), .b(new_n189_), .O(new_n283_));
  AND      g267(.a(new_n283_), .b(i_2_2_63_0), .O(new_n284_));
  NAND     g268(.a(new_n132_), .b(i_2_2_129_0), .O(new_n285_));
  NAND     g269(.a(new_n285_), .b(new_n60_), .O(new_n286_));
  AND      g270(.a(new_n286_), .b(i_2_2_91_0), .O(new_n287_));
  AND      g271(.a(new_n19_), .b(i_2_2_129_0), .O(new_n288_));
  OR       g272(.a(new_n288_), .b(i_2_2_134_0), .O(new_n289_));
  OR       g273(.a(i_2_2_134_0), .b(i_2_2_116_0), .O(new_n290_));
  AND      g274(.a(new_n290_), .b(new_n19_), .O(new_n291_));
  OR       g275(.a(new_n291_), .b(new_n21_), .O(new_n292_));
  AND      g276(.a(new_n292_), .b(new_n289_), .O(new_n293_));
  OR       g277(.a(new_n293_), .b(new_n287_), .O(new_n294_));
  OR       g278(.a(new_n294_), .b(new_n284_), .O(new_n295_));
  AND      g279(.a(new_n295_), .b(i_2_2_137_0), .O(new_n296_));
  AND      g280(.a(new_n209_), .b(new_n132_), .O(new_n297_));
  AND      g281(.a(new_n297_), .b(new_n200_), .O(new_n298_));
  NAND     g282(.a(new_n132_), .b(new_n67_), .O(new_n299_));
  NOT      g283(.a(new_n42_), .O(new_n300_));
  AND      g284(.a(new_n158_), .b(new_n300_), .O(new_n301_));
  OR       g285(.a(new_n301_), .b(new_n166_), .O(new_n302_));
  NAND     g286(.a(new_n302_), .b(new_n299_), .O(new_n303_));
  AND      g287(.a(new_n303_), .b(i_2_2_63_0), .O(new_n304_));
  OR       g288(.a(new_n189_), .b(new_n39_), .O(new_n305_));
  NOT      g289(.a(new_n159_), .O(new_n306_));
  OR       g290(.a(new_n306_), .b(new_n91_), .O(new_n307_));
  AND      g291(.a(new_n307_), .b(i_2_2_116_0), .O(new_n308_));
  AND      g292(.a(new_n308_), .b(new_n305_), .O(new_n309_));
  OR       g293(.a(new_n309_), .b(new_n304_), .O(new_n310_));
  AND      g294(.a(new_n310_), .b(new_n19_), .O(new_n311_));
  OR       g295(.a(new_n311_), .b(new_n298_), .O(new_n312_));
  OR       g296(.a(new_n312_), .b(new_n296_), .O(new_n313_));
  AND      g297(.a(new_n313_), .b(i_2_2_58_0), .O(new_n314_));
  OR       g298(.a(new_n173_), .b(new_n19_), .O(new_n315_));
  AND      g299(.a(new_n315_), .b(new_n172_), .O(new_n316_));
  NOT      g300(.a(new_n227_), .O(new_n317_));
  NAND     g301(.a(i_2_2_147_0), .b(i_2_2_63_0), .O(new_n318_));
  AND      g302(.a(new_n318_), .b(i_2_2_107_0), .O(new_n319_));
  OR       g303(.a(new_n49_), .b(i_2_2_116_0), .O(new_n320_));
  OR       g304(.a(new_n320_), .b(new_n319_), .O(new_n321_));
  NAND     g305(.a(new_n321_), .b(new_n317_), .O(new_n322_));
  OR       g306(.a(new_n322_), .b(new_n316_), .O(new_n323_));
  AND      g307(.a(new_n323_), .b(i_2_2_91_0), .O(new_n324_));
  NAND     g308(.a(i_2_2_129_0), .b(i_2_2_63_0), .O(new_n325_));
  NAND     g309(.a(new_n325_), .b(i_2_2_147_0), .O(new_n326_));
  OR       g310(.a(new_n173_), .b(new_n189_), .O(new_n327_));
  AND      g311(.a(new_n327_), .b(new_n326_), .O(new_n328_));
  AND      g312(.a(new_n288_), .b(i_2_2_63_0), .O(new_n329_));
  OR       g313(.a(i_2_2_134_0), .b(i_2_2_58_0), .O(new_n330_));
  OR       g314(.a(new_n330_), .b(new_n329_), .O(new_n331_));
  OR       g315(.a(new_n331_), .b(new_n328_), .O(new_n332_));
  AND      g316(.a(new_n332_), .b(i_2_2_116_0), .O(new_n333_));
  AND      g317(.a(new_n227_), .b(i_2_2_63_0), .O(new_n334_));
  AND      g318(.a(new_n326_), .b(i_2_2_58_0), .O(new_n335_));
  OR       g319(.a(new_n148_), .b(new_n19_), .O(new_n336_));
  AND      g320(.a(new_n336_), .b(i_2_2_134_0), .O(new_n337_));
  OR       g321(.a(new_n337_), .b(new_n335_), .O(new_n338_));
  AND      g322(.a(new_n338_), .b(new_n21_), .O(new_n339_));
  OR       g323(.a(new_n339_), .b(new_n334_), .O(new_n340_));
  OR       g324(.a(new_n340_), .b(new_n333_), .O(new_n341_));
  OR       g325(.a(new_n341_), .b(new_n324_), .O(new_n342_));
  AND      g326(.a(new_n342_), .b(new_n39_), .O(new_n343_));
  AND      g327(.a(new_n19_), .b(i_2_2_139_0), .O(new_n344_));
  NAND     g328(.a(new_n344_), .b(i_2_2_58_0), .O(new_n345_));
  NAND     g329(.a(new_n345_), .b(new_n56_), .O(new_n346_));
  AND      g330(.a(new_n346_), .b(new_n115_), .O(new_n347_));
  NOT      g331(.a(new_n288_), .O(new_n348_));
  OR       g332(.a(new_n348_), .b(new_n174_), .O(new_n349_));
  AND      g333(.a(i_2_2_134_0), .b(i_2_2_116_0), .O(new_n350_));
  NAND     g334(.a(new_n350_), .b(new_n315_), .O(new_n351_));
  NAND     g335(.a(new_n351_), .b(new_n349_), .O(new_n352_));
  OR       g336(.a(new_n352_), .b(new_n347_), .O(new_n353_));
  OR       g337(.a(new_n353_), .b(new_n343_), .O(new_n354_));
  AND      g338(.a(new_n354_), .b(i_2_2_137_0), .O(new_n355_));
  OR       g339(.a(new_n355_), .b(new_n314_), .O(new_n356_));
  AND      g340(.a(new_n356_), .b(new_n20_), .O(new_n357_));
  AND      g341(.a(i_2_2_137_0), .b(i_2_2_58_0), .O(new_n358_));
  AND      g342(.a(new_n180_), .b(new_n60_), .O(new_n359_));
  AND      g343(.a(i_2_2_116_0), .b(i_2_2_63_0), .O(new_n360_));
  AND      g344(.a(new_n360_), .b(new_n177_), .O(new_n361_));
  OR       g345(.a(new_n361_), .b(new_n359_), .O(new_n362_));
  AND      g346(.a(new_n362_), .b(new_n358_), .O(new_n363_));
  AND      g347(.a(i_2_2_116_0), .b(i_2_2_58_0), .O(new_n364_));
  OR       g348(.a(new_n140_), .b(new_n23_), .O(new_n365_));
  AND      g349(.a(new_n365_), .b(new_n364_), .O(new_n366_));
  AND      g350(.a(new_n202_), .b(i_2_2_58_0), .O(new_n367_));
  OR       g351(.a(new_n364_), .b(new_n149_), .O(new_n368_));
  OR       g352(.a(new_n368_), .b(new_n367_), .O(new_n369_));
  AND      g353(.a(new_n369_), .b(new_n19_), .O(new_n370_));
  OR       g354(.a(new_n370_), .b(new_n366_), .O(new_n371_));
  AND      g355(.a(new_n371_), .b(i_2_2_134_0), .O(new_n372_));
  AND      g356(.a(new_n147_), .b(i_2_2_129_0), .O(new_n373_));
  AND      g357(.a(new_n373_), .b(new_n358_), .O(new_n374_));
  OR       g358(.a(new_n373_), .b(new_n233_), .O(new_n375_));
  AND      g359(.a(new_n375_), .b(i_2_2_139_0), .O(new_n376_));
  AND      g360(.a(new_n274_), .b(new_n264_), .O(new_n377_));
  OR       g361(.a(new_n377_), .b(new_n258_), .O(new_n378_));
  OR       g362(.a(new_n378_), .b(new_n376_), .O(new_n379_));
  AND      g363(.a(new_n379_), .b(i_2_2_58_0), .O(new_n380_));
  AND      g364(.a(new_n260_), .b(new_n147_), .O(new_n381_));
  AND      g365(.a(new_n381_), .b(new_n140_), .O(new_n382_));
  OR       g366(.a(new_n382_), .b(new_n380_), .O(new_n383_));
  AND      g367(.a(new_n383_), .b(new_n19_), .O(new_n384_));
  OR       g368(.a(new_n384_), .b(new_n374_), .O(new_n385_));
  OR       g369(.a(new_n385_), .b(new_n372_), .O(new_n386_));
  AND      g370(.a(new_n386_), .b(new_n21_), .O(new_n387_));
  OR       g371(.a(new_n387_), .b(new_n363_), .O(new_n388_));
  AND      g372(.a(new_n388_), .b(new_n39_), .O(new_n389_));
  OR       g373(.a(new_n389_), .b(new_n357_), .O(new_n390_));
  OR       g374(.a(new_n390_), .b(new_n278_), .O(new_n391_));
  AND      g375(.a(new_n391_), .b(new_n18_), .O(new_n392_));
  AND      g376(.a(i_2_2_134_0), .b(i_2_2_91_0), .O(new_n393_));
  AND      g377(.a(i_2_2_129_0), .b(new_n20_), .O(new_n394_));
  OR       g378(.a(new_n394_), .b(new_n393_), .O(new_n395_));
  AND      g379(.a(new_n395_), .b(new_n257_), .O(new_n396_));
  OR       g380(.a(i_2_2_147_0), .b(new_n40_), .O(new_n397_));
  OR       g381(.a(new_n19_), .b(i_2_2_82_0), .O(new_n398_));
  NAND     g382(.a(new_n398_), .b(new_n397_), .O(new_n399_));
  AND      g383(.a(new_n399_), .b(new_n20_), .O(new_n400_));
  OR       g384(.a(new_n19_), .b(i_2_2_91_0), .O(new_n401_));
  AND      g385(.a(new_n401_), .b(new_n152_), .O(new_n402_));
  OR       g386(.a(new_n402_), .b(new_n400_), .O(new_n403_));
  AND      g387(.a(new_n403_), .b(i_2_2_139_0), .O(new_n404_));
  OR       g388(.a(i_2_2_139_0), .b(i_2_2_82_0), .O(new_n405_));
  AND      g389(.a(new_n405_), .b(i_2_2_60_0), .O(new_n406_));
  OR       g390(.a(new_n406_), .b(new_n397_), .O(new_n407_));
  NAND     g391(.a(new_n407_), .b(new_n61_), .O(new_n408_));
  AND      g392(.a(new_n408_), .b(i_2_2_129_0), .O(new_n409_));
  AND      g393(.a(new_n19_), .b(i_2_2_134_0), .O(new_n410_));
  AND      g394(.a(new_n410_), .b(new_n20_), .O(new_n411_));
  OR       g395(.a(new_n411_), .b(new_n409_), .O(new_n412_));
  OR       g396(.a(new_n412_), .b(new_n404_), .O(new_n413_));
  AND      g397(.a(new_n413_), .b(i_2_2_63_0), .O(new_n414_));
  OR       g398(.a(new_n414_), .b(new_n396_), .O(new_n415_));
  AND      g399(.a(new_n415_), .b(new_n21_), .O(new_n416_));
  OR       g400(.a(new_n257_), .b(new_n180_), .O(new_n417_));
  AND      g401(.a(i_2_2_147_0), .b(new_n39_), .O(new_n418_));
  OR       g402(.a(new_n410_), .b(new_n418_), .O(new_n419_));
  AND      g403(.a(new_n419_), .b(new_n20_), .O(new_n420_));
  AND      g404(.a(new_n420_), .b(new_n417_), .O(new_n421_));
  AND      g405(.a(i_2_2_139_0), .b(new_n39_), .O(new_n422_));
  AND      g406(.a(new_n422_), .b(i_2_2_91_0), .O(new_n423_));
  NAND     g407(.a(new_n288_), .b(i_2_2_134_0), .O(new_n424_));
  NOT      g408(.a(new_n424_), .O(new_n425_));
  AND      g409(.a(new_n425_), .b(new_n423_), .O(new_n426_));
  OR       g410(.a(new_n426_), .b(new_n421_), .O(new_n427_));
  OR       g411(.a(new_n427_), .b(new_n416_), .O(new_n428_));
  AND      g412(.a(new_n428_), .b(i_2_2_116_0), .O(new_n429_));
  NOT      g413(.a(new_n49_), .O(new_n430_));
  OR       g414(.a(i_2_2_91_0), .b(i_2_2_82_0), .O(new_n431_));
  AND      g415(.a(new_n431_), .b(new_n430_), .O(new_n432_));
  AND      g416(.a(new_n422_), .b(new_n274_), .O(new_n433_));
  OR       g417(.a(new_n433_), .b(new_n432_), .O(new_n434_));
  AND      g418(.a(new_n411_), .b(new_n21_), .O(new_n435_));
  AND      g419(.a(new_n435_), .b(new_n434_), .O(new_n436_));
  OR       g420(.a(new_n436_), .b(new_n429_), .O(new_n437_));
  AND      g421(.a(new_n437_), .b(i_2_2_137_0), .O(new_n438_));
  OR       g422(.a(new_n344_), .b(new_n39_), .O(new_n439_));
  OR       g423(.a(new_n439_), .b(new_n393_), .O(new_n440_));
  AND      g424(.a(new_n440_), .b(i_2_2_137_0), .O(new_n441_));
  AND      g425(.a(new_n19_), .b(i_2_2_91_0), .O(new_n442_));
  AND      g426(.a(new_n442_), .b(i_2_2_139_0), .O(new_n443_));
  AND      g427(.a(new_n443_), .b(i_2_2_134_0), .O(new_n444_));
  OR       g428(.a(new_n444_), .b(new_n441_), .O(new_n445_));
  AND      g429(.a(new_n445_), .b(i_2_2_129_0), .O(new_n446_));
  AND      g430(.a(new_n257_), .b(new_n22_), .O(new_n447_));
  OR       g431(.a(new_n447_), .b(new_n119_), .O(new_n448_));
  OR       g432(.a(new_n448_), .b(new_n446_), .O(new_n449_));
  AND      g433(.a(new_n449_), .b(i_2_2_63_0), .O(new_n450_));
  AND      g434(.a(new_n238_), .b(i_2_2_134_0), .O(new_n451_));
  OR       g435(.a(i_2_2_139_0), .b(i_2_2_134_0), .O(new_n452_));
  AND      g436(.a(new_n452_), .b(new_n91_), .O(new_n453_));
  OR       g437(.a(new_n453_), .b(new_n260_), .O(new_n454_));
  AND      g438(.a(new_n454_), .b(new_n39_), .O(new_n455_));
  OR       g439(.a(new_n455_), .b(new_n451_), .O(new_n456_));
  OR       g440(.a(new_n456_), .b(new_n450_), .O(new_n457_));
  AND      g441(.a(new_n457_), .b(new_n20_), .O(new_n458_));
  OR       g442(.a(new_n397_), .b(new_n62_), .O(new_n459_));
  NAND     g443(.a(new_n459_), .b(new_n41_), .O(new_n460_));
  AND      g444(.a(new_n460_), .b(new_n39_), .O(new_n461_));
  AND      g445(.a(new_n238_), .b(i_2_2_91_0), .O(new_n462_));
  OR       g446(.a(new_n462_), .b(new_n461_), .O(new_n463_));
  AND      g447(.a(new_n463_), .b(i_2_2_129_0), .O(new_n464_));
  NOT      g448(.a(new_n405_), .O(new_n465_));
  AND      g449(.a(new_n19_), .b(i_2_2_63_0), .O(new_n466_));
  AND      g450(.a(new_n466_), .b(i_2_2_139_0), .O(new_n467_));
  OR       g451(.a(new_n467_), .b(new_n465_), .O(new_n468_));
  AND      g452(.a(new_n468_), .b(i_2_2_137_0), .O(new_n469_));
  OR       g453(.a(new_n469_), .b(new_n464_), .O(new_n470_));
  AND      g454(.a(new_n470_), .b(i_2_2_134_0), .O(new_n471_));
  AND      g455(.a(i_2_2_137_0), .b(new_n115_), .O(new_n472_));
  AND      g456(.a(new_n472_), .b(new_n91_), .O(new_n473_));
  AND      g457(.a(new_n473_), .b(new_n257_), .O(new_n474_));
  OR       g458(.a(new_n474_), .b(new_n471_), .O(new_n475_));
  OR       g459(.a(new_n475_), .b(new_n458_), .O(new_n476_));
  AND      g460(.a(new_n476_), .b(i_2_2_116_0), .O(new_n477_));
  AND      g461(.a(new_n91_), .b(i_2_2_147_0), .O(new_n478_));
  OR       g462(.a(new_n394_), .b(i_2_2_139_0), .O(new_n479_));
  AND      g463(.a(new_n479_), .b(new_n478_), .O(new_n480_));
  OR       g464(.a(new_n480_), .b(new_n99_), .O(new_n481_));
  AND      g465(.a(new_n481_), .b(i_2_2_116_0), .O(new_n482_));
  OR       g466(.a(new_n442_), .b(i_2_2_116_0), .O(new_n483_));
  AND      g467(.a(new_n483_), .b(new_n325_), .O(new_n484_));
  NAND     g468(.a(new_n459_), .b(new_n98_), .O(new_n485_));
  OR       g469(.a(new_n485_), .b(new_n484_), .O(new_n486_));
  AND      g470(.a(new_n486_), .b(i_2_2_137_0), .O(new_n487_));
  OR       g471(.a(new_n487_), .b(new_n482_), .O(new_n488_));
  AND      g472(.a(new_n488_), .b(i_2_2_134_0), .O(new_n489_));
  AND      g473(.a(i_2_2_137_0), .b(new_n20_), .O(new_n490_));
  OR       g474(.a(new_n19_), .b(i_2_2_139_0), .O(new_n491_));
  AND      g475(.a(new_n491_), .b(i_2_2_116_0), .O(new_n492_));
  OR       g476(.a(new_n492_), .b(new_n423_), .O(new_n493_));
  AND      g477(.a(new_n493_), .b(new_n490_), .O(new_n494_));
  OR       g478(.a(new_n494_), .b(new_n489_), .O(new_n495_));
  AND      g479(.a(new_n495_), .b(new_n21_), .O(new_n496_));
  AND      g480(.a(new_n460_), .b(new_n20_), .O(new_n497_));
  AND      g481(.a(new_n442_), .b(new_n233_), .O(new_n498_));
  OR       g482(.a(new_n498_), .b(new_n497_), .O(new_n499_));
  AND      g483(.a(new_n152_), .b(i_2_2_129_0), .O(new_n500_));
  AND      g484(.a(new_n500_), .b(new_n499_), .O(new_n501_));
  OR       g485(.a(new_n501_), .b(new_n496_), .O(new_n502_));
  OR       g486(.a(new_n502_), .b(new_n477_), .O(new_n503_));
  AND      g487(.a(new_n503_), .b(i_2_2_58_0), .O(new_n504_));
  OR       g488(.a(i_2_2_108_0), .b(i_2_2_91_0), .O(new_n505_));
  AND      g489(.a(new_n505_), .b(new_n62_), .O(new_n506_));
  OR       g490(.a(new_n506_), .b(new_n20_), .O(new_n507_));
  AND      g491(.a(new_n425_), .b(new_n297_), .O(new_n508_));
  AND      g492(.a(new_n508_), .b(new_n507_), .O(new_n509_));
  OR       g493(.a(new_n509_), .b(new_n504_), .O(new_n510_));
  OR       g494(.a(new_n510_), .b(new_n438_), .O(new_n511_));
  OR       g495(.a(new_n511_), .b(new_n392_), .O(new_n512_));
  AND      g496(.a(new_n512_), .b(new_n157_), .O(new_n513_));
  AND      g497(.a(new_n44_), .b(i_2_2_107_0), .O(new_n514_));
  AND      g498(.a(new_n514_), .b(new_n109_), .O(new_n515_));
  NAND     g499(.a(new_n274_), .b(i_2_2_116_0), .O(new_n516_));
  NAND     g500(.a(i_2_2_129_0), .b(i_2_2_108_0), .O(new_n517_));
  OR       g501(.a(new_n517_), .b(new_n290_), .O(new_n518_));
  NAND     g502(.a(new_n518_), .b(new_n516_), .O(new_n519_));
  OR       g503(.a(i_2_2_147_0), .b(i_2_2_107_0), .O(new_n520_));
  NOT      g504(.a(new_n520_), .O(new_n521_));
  AND      g505(.a(new_n521_), .b(new_n519_), .O(new_n522_));
  OR       g506(.a(new_n522_), .b(new_n515_), .O(new_n523_));
  AND      g507(.a(new_n523_), .b(i_2_2_137_0), .O(new_n524_));
  AND      g508(.a(i_2_2_108_0), .b(i_2_2_107_0), .O(new_n525_));
  AND      g509(.a(new_n525_), .b(new_n41_), .O(new_n526_));
  OR       g510(.a(new_n526_), .b(new_n238_), .O(new_n527_));
  AND      g511(.a(new_n147_), .b(new_n44_), .O(new_n528_));
  AND      g512(.a(new_n528_), .b(new_n527_), .O(new_n529_));
  OR       g513(.a(new_n529_), .b(new_n524_), .O(new_n530_));
  AND      g514(.a(new_n530_), .b(i_2_2_58_0), .O(new_n531_));
  OR       g515(.a(new_n177_), .b(new_n108_), .O(new_n532_));
  NOT      g516(.a(new_n532_), .O(new_n533_));
  AND      g517(.a(new_n466_), .b(i_2_2_108_0), .O(new_n534_));
  OR       g518(.a(i_2_2_137_0), .b(i_2_2_107_0), .O(new_n535_));
  NOT      g519(.a(new_n535_), .O(new_n536_));
  AND      g520(.a(new_n536_), .b(new_n44_), .O(new_n537_));
  AND      g521(.a(new_n537_), .b(new_n534_), .O(new_n538_));
  AND      g522(.a(new_n538_), .b(new_n533_), .O(new_n539_));
  OR       g523(.a(new_n539_), .b(new_n531_), .O(new_n540_));
  AND      g524(.a(new_n540_), .b(new_n20_), .O(new_n541_));
  NOT      g525(.a(new_n452_), .O(new_n542_));
  AND      g526(.a(new_n542_), .b(new_n258_), .O(new_n543_));
  AND      g527(.a(new_n543_), .b(new_n55_), .O(new_n544_));
  AND      g528(.a(new_n544_), .b(new_n534_), .O(new_n545_));
  OR       g529(.a(new_n545_), .b(new_n541_), .O(new_n546_));
  AND      g530(.a(new_n546_), .b(new_n39_), .O(new_n547_));
  AND      g531(.a(i_2_2_63_0), .b(i_2_2_58_0), .O(new_n548_));
  AND      g532(.a(new_n91_), .b(new_n20_), .O(new_n549_));
  AND      g533(.a(new_n549_), .b(new_n548_), .O(new_n550_));
  NOT      g534(.a(new_n247_), .O(new_n551_));
  OR       g535(.a(new_n551_), .b(new_n132_), .O(new_n552_));
  OR       g536(.a(new_n525_), .b(i_2_2_147_0), .O(new_n553_));
  AND      g537(.a(new_n553_), .b(new_n119_), .O(new_n554_));
  AND      g538(.a(new_n554_), .b(new_n552_), .O(new_n555_));
  AND      g539(.a(new_n555_), .b(new_n550_), .O(new_n556_));
  OR       g540(.a(new_n556_), .b(new_n547_), .O(new_n557_));
  OR       g541(.a(new_n557_), .b(new_n513_), .O(new_n558_));
  OR       g542(.a(new_n558_), .b(new_n156_), .O(new_n559_));
  AND      g543(.a(new_n559_), .b(new_n17_), .O(new_n560_));
  OR       g544(.a(i_2_2_147_0), .b(i_2_2_60_0), .O(new_n561_));
  NOT      g545(.a(new_n561_), .O(new_n562_));
  OR       g546(.a(new_n264_), .b(new_n212_), .O(new_n563_));
  OR       g547(.a(new_n158_), .b(i_2_2_82_0), .O(new_n564_));
  NAND     g548(.a(new_n564_), .b(new_n563_), .O(new_n565_));
  AND      g549(.a(new_n565_), .b(new_n562_), .O(new_n566_));
  NOT      g550(.a(new_n264_), .O(new_n567_));
  AND      g551(.a(new_n567_), .b(i_2_2_147_0), .O(new_n568_));
  AND      g552(.a(new_n568_), .b(new_n423_), .O(new_n569_));
  OR       g553(.a(new_n569_), .b(new_n566_), .O(new_n570_));
  AND      g554(.a(new_n570_), .b(i_2_2_129_0), .O(new_n571_));
  AND      g555(.a(i_2_2_147_0), .b(new_n48_), .O(new_n572_));
  AND      g556(.a(new_n572_), .b(new_n99_), .O(new_n573_));
  AND      g557(.a(new_n573_), .b(new_n138_), .O(new_n574_));
  OR       g558(.a(new_n574_), .b(new_n571_), .O(new_n575_));
  AND      g559(.a(new_n575_), .b(new_n21_), .O(new_n576_));
  AND      g560(.a(new_n23_), .b(i_2_2_147_0), .O(new_n577_));
  AND      g561(.a(new_n109_), .b(new_n99_), .O(new_n578_));
  AND      g562(.a(new_n578_), .b(new_n577_), .O(new_n579_));
  OR       g563(.a(new_n579_), .b(new_n576_), .O(new_n580_));
  AND      g564(.a(new_n580_), .b(new_n548_), .O(new_n581_));
  OR       g565(.a(new_n348_), .b(new_n194_), .O(new_n582_));
  NAND     g566(.a(new_n582_), .b(new_n98_), .O(new_n583_));
  AND      g567(.a(new_n583_), .b(i_2_2_63_0), .O(new_n584_));
  AND      g568(.a(new_n491_), .b(new_n20_), .O(new_n585_));
  AND      g569(.a(new_n344_), .b(new_n40_), .O(new_n586_));
  OR       g570(.a(new_n586_), .b(new_n585_), .O(new_n587_));
  AND      g571(.a(new_n587_), .b(new_n39_), .O(new_n588_));
  OR       g572(.a(new_n588_), .b(new_n584_), .O(new_n589_));
  AND      g573(.a(new_n589_), .b(i_2_2_58_0), .O(new_n590_));
  AND      g574(.a(new_n72_), .b(i_2_2_129_0), .O(new_n591_));
  OR       g575(.a(new_n591_), .b(new_n21_), .O(new_n592_));
  NAND     g576(.a(new_n42_), .b(new_n21_), .O(new_n593_));
  AND      g577(.a(i_2_2_147_0), .b(i_2_2_60_0), .O(new_n594_));
  AND      g578(.a(new_n594_), .b(new_n593_), .O(new_n595_));
  AND      g579(.a(new_n595_), .b(new_n592_), .O(new_n596_));
  OR       g580(.a(new_n596_), .b(new_n590_), .O(new_n597_));
  AND      g581(.a(new_n597_), .b(i_2_2_116_0), .O(new_n598_));
  AND      g582(.a(new_n573_), .b(new_n109_), .O(new_n599_));
  NOT      g583(.a(new_n478_), .O(new_n600_));
  OR       g584(.a(new_n600_), .b(new_n243_), .O(new_n601_));
  NAND     g585(.a(new_n601_), .b(new_n561_), .O(new_n602_));
  AND      g586(.a(i_2_2_139_0), .b(i_2_2_58_0), .O(new_n603_));
  AND      g587(.a(new_n603_), .b(new_n602_), .O(new_n604_));
  OR       g588(.a(new_n604_), .b(new_n599_), .O(new_n605_));
  AND      g589(.a(new_n605_), .b(new_n21_), .O(new_n606_));
  NOT      g590(.a(new_n243_), .O(new_n607_));
  AND      g591(.a(new_n467_), .b(new_n607_), .O(new_n608_));
  AND      g592(.a(new_n608_), .b(new_n591_), .O(new_n609_));
  OR       g593(.a(new_n609_), .b(new_n606_), .O(new_n610_));
  OR       g594(.a(new_n610_), .b(new_n598_), .O(new_n611_));
  AND      g595(.a(new_n611_), .b(i_2_2_137_0), .O(new_n612_));
  OR       g596(.a(new_n612_), .b(new_n581_), .O(new_n613_));
  AND      g597(.a(new_n613_), .b(new_n157_), .O(new_n614_));
  OR       g598(.a(new_n279_), .b(new_n246_), .O(new_n615_));
  OR       g599(.a(new_n397_), .b(i_2_2_58_0), .O(new_n616_));
  OR       g600(.a(new_n616_), .b(new_n285_), .O(new_n617_));
  NAND     g601(.a(new_n617_), .b(new_n615_), .O(new_n618_));
  AND      g602(.a(new_n490_), .b(new_n148_), .O(new_n619_));
  AND      g603(.a(new_n619_), .b(new_n618_), .O(new_n620_));
  OR       g604(.a(new_n620_), .b(new_n614_), .O(new_n621_));
  AND      g605(.a(new_n621_), .b(i_2_2_134_0), .O(new_n622_));
  AND      g606(.a(new_n577_), .b(new_n85_), .O(new_n623_));
  AND      g607(.a(new_n227_), .b(new_n209_), .O(new_n624_));
  AND      g608(.a(new_n624_), .b(new_n479_), .O(new_n625_));
  OR       g609(.a(new_n625_), .b(new_n623_), .O(new_n626_));
  NOT      g610(.a(new_n94_), .O(new_n627_));
  AND      g611(.a(new_n258_), .b(new_n157_), .O(new_n628_));
  AND      g612(.a(new_n628_), .b(new_n627_), .O(new_n629_));
  AND      g613(.a(new_n629_), .b(new_n626_), .O(new_n630_));
  OR       g614(.a(new_n630_), .b(new_n622_), .O(new_n631_));
  AND      g615(.a(new_n631_), .b(new_n18_), .O(new_n632_));
  NAND     g616(.a(new_n490_), .b(i_2_2_91_0), .O(new_n633_));
  AND      g617(.a(new_n178_), .b(new_n108_), .O(new_n634_));
  AND      g618(.a(new_n532_), .b(i_2_2_60_0), .O(new_n635_));
  OR       g619(.a(new_n635_), .b(new_n60_), .O(new_n636_));
  OR       g620(.a(new_n636_), .b(new_n634_), .O(new_n637_));
  NAND     g621(.a(new_n637_), .b(new_n633_), .O(new_n638_));
  AND      g622(.a(new_n638_), .b(new_n17_), .O(new_n639_));
  AND      g623(.a(new_n490_), .b(i_2_2_139_0), .O(new_n640_));
  AND      g624(.a(new_n640_), .b(new_n607_), .O(new_n641_));
  OR       g625(.a(new_n641_), .b(new_n639_), .O(new_n642_));
  AND      g626(.a(new_n642_), .b(new_n19_), .O(new_n643_));
  NAND     g627(.a(i_2_2_137_0), .b(i_2_2_108_0), .O(new_n644_));
  OR       g628(.a(new_n644_), .b(new_n600_), .O(new_n645_));
  OR       g629(.a(new_n108_), .b(i_2_2_113_0), .O(new_n646_));
  OR       g630(.a(i_2_2_147_0), .b(i_2_2_91_0), .O(new_n647_));
  OR       g631(.a(new_n647_), .b(new_n646_), .O(new_n648_));
  NAND     g632(.a(new_n648_), .b(new_n645_), .O(new_n649_));
  AND      g633(.a(new_n649_), .b(i_2_2_60_0), .O(new_n650_));
  OR       g634(.a(new_n451_), .b(new_n411_), .O(new_n651_));
  AND      g635(.a(new_n490_), .b(i_2_2_116_0), .O(new_n652_));
  OR       g636(.a(new_n652_), .b(new_n17_), .O(new_n653_));
  AND      g637(.a(new_n653_), .b(new_n651_), .O(new_n654_));
  OR       g638(.a(new_n654_), .b(new_n650_), .O(new_n655_));
  AND      g639(.a(new_n655_), .b(i_2_2_139_0), .O(new_n656_));
  AND      g640(.a(new_n561_), .b(new_n75_), .O(new_n657_));
  OR       g641(.a(new_n657_), .b(new_n646_), .O(new_n658_));
  NOT      g642(.a(new_n572_), .O(new_n659_));
  AND      g643(.a(new_n659_), .b(new_n424_), .O(new_n660_));
  NAND     g644(.a(new_n124_), .b(new_n49_), .O(new_n661_));
  NAND     g645(.a(new_n490_), .b(new_n661_), .O(new_n662_));
  OR       g646(.a(new_n662_), .b(new_n660_), .O(new_n663_));
  NAND     g647(.a(new_n663_), .b(new_n658_), .O(new_n664_));
  AND      g648(.a(new_n664_), .b(i_2_2_91_0), .O(new_n665_));
  AND      g649(.a(new_n290_), .b(new_n20_), .O(new_n666_));
  OR       g650(.a(new_n666_), .b(new_n27_), .O(new_n667_));
  AND      g651(.a(new_n288_), .b(new_n17_), .O(new_n668_));
  AND      g652(.a(new_n668_), .b(new_n667_), .O(new_n669_));
  OR       g653(.a(new_n669_), .b(new_n665_), .O(new_n670_));
  OR       g654(.a(new_n670_), .b(new_n656_), .O(new_n671_));
  AND      g655(.a(new_n671_), .b(new_n39_), .O(new_n672_));
  OR       g656(.a(new_n672_), .b(new_n643_), .O(new_n673_));
  AND      g657(.a(new_n673_), .b(i_2_2_63_0), .O(new_n674_));
  NOT      g658(.a(new_n645_), .O(new_n675_));
  AND      g659(.a(i_2_2_82_0), .b(new_n20_), .O(new_n676_));
  AND      g660(.a(new_n676_), .b(new_n44_), .O(new_n677_));
  AND      g661(.a(new_n677_), .b(new_n675_), .O(new_n678_));
  OR       g662(.a(new_n678_), .b(new_n674_), .O(new_n679_));
  AND      g663(.a(new_n679_), .b(new_n21_), .O(new_n680_));
  AND      g664(.a(new_n562_), .b(new_n422_), .O(new_n681_));
  AND      g665(.a(new_n681_), .b(new_n126_), .O(new_n682_));
  OR       g666(.a(new_n682_), .b(new_n680_), .O(new_n683_));
  AND      g667(.a(i_2_2_58_0), .b(new_n157_), .O(new_n684_));
  AND      g668(.a(new_n684_), .b(new_n683_), .O(new_n685_));
  OR       g669(.a(new_n685_), .b(new_n632_), .O(new_n686_));
  OR       g670(.a(new_n686_), .b(new_n560_), .O(o_2_2_0_0));
endmodule


