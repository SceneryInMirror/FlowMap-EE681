module kernel_2_6 ( 
    i_2_6_5_0, i_2_6_32_0, i_2_6_33_0, i_2_6_34_0, i_2_6_40_0, i_2_6_51_0,
    i_2_6_62_0, i_2_6_63_0, i_2_6_84_0, i_2_6_110_0, i_2_6_111_0,
    i_2_6_118_0, i_2_6_120_0, i_2_6_124_0, i_2_6_142_0,
    o_2_6_0_0  );
  input  i_2_6_5_0, i_2_6_32_0, i_2_6_33_0, i_2_6_34_0, i_2_6_40_0,
    i_2_6_51_0, i_2_6_62_0, i_2_6_63_0, i_2_6_84_0, i_2_6_110_0,
    i_2_6_111_0, i_2_6_118_0, i_2_6_120_0, i_2_6_124_0, i_2_6_142_0;
  output o_2_6_0_0;
  assign o_2_6_0_0 = (~i_2_6_120_0 & ((i_2_6_5_0 & ((~i_2_6_51_0 & ((i_2_6_33_0 & ((i_2_6_62_0 & ((i_2_6_34_0 & ((i_2_6_40_0 & ((~i_2_6_118_0 & ~i_2_6_124_0) | (~i_2_6_84_0 & i_2_6_142_0))) | (i_2_6_111_0 & (i_2_6_63_0 | (i_2_6_32_0 & ~i_2_6_40_0 & i_2_6_110_0))) | (~i_2_6_40_0 & (((i_2_6_32_0 | i_2_6_63_0) & (~i_2_6_84_0 | ~i_2_6_118_0)) | (i_2_6_32_0 & i_2_6_63_0))) | (i_2_6_63_0 & ((i_2_6_32_0 & (~i_2_6_124_0 | i_2_6_142_0)) | (~i_2_6_84_0 & i_2_6_110_0))) | (~i_2_6_124_0 & ((i_2_6_110_0 & (~i_2_6_118_0 | i_2_6_142_0)) | (~i_2_6_118_0 & i_2_6_142_0))))) | (i_2_6_110_0 & ((~i_2_6_118_0 & ((i_2_6_32_0 & ((~i_2_6_63_0 & ~i_2_6_111_0 & i_2_6_124_0) | (~i_2_6_40_0 & i_2_6_63_0 & ~i_2_6_124_0))) | ~i_2_6_84_0 | (~i_2_6_63_0 & i_2_6_124_0 & i_2_6_142_0))) | (i_2_6_63_0 & ((~i_2_6_40_0 & ~i_2_6_124_0 & (~i_2_6_84_0 | i_2_6_111_0)) | (i_2_6_32_0 & ~i_2_6_84_0 & i_2_6_111_0))))) | (i_2_6_111_0 & ((~i_2_6_118_0 & ((~i_2_6_84_0 & i_2_6_124_0) | (i_2_6_32_0 & i_2_6_63_0 & ~i_2_6_124_0))) | (i_2_6_63_0 & ((i_2_6_32_0 & ~i_2_6_84_0 & (~i_2_6_40_0 | ~i_2_6_124_0)) | (i_2_6_118_0 & ~i_2_6_124_0 & i_2_6_142_0))) | (~i_2_6_40_0 & i_2_6_142_0 & ((i_2_6_84_0 & ~i_2_6_110_0 & i_2_6_124_0) | (~i_2_6_84_0 & ~i_2_6_124_0))))) | (i_2_6_32_0 & ~i_2_6_40_0 & i_2_6_63_0 & ~i_2_6_118_0 & ~i_2_6_124_0 & i_2_6_142_0))) | (~i_2_6_118_0 & ((i_2_6_34_0 & (i_2_6_111_0 | (i_2_6_32_0 & i_2_6_63_0))) | (~i_2_6_111_0 & ((~i_2_6_32_0 & i_2_6_40_0 & i_2_6_110_0) | (~i_2_6_124_0 & i_2_6_142_0 & ~i_2_6_84_0 & ~i_2_6_110_0))) | (i_2_6_32_0 & ((i_2_6_63_0 & ((~i_2_6_40_0 & (~i_2_6_84_0 | (i_2_6_111_0 & ~i_2_6_142_0))) | (~i_2_6_84_0 & ~i_2_6_124_0) | (i_2_6_111_0 & ((~i_2_6_124_0 & i_2_6_142_0) | (i_2_6_110_0 & i_2_6_124_0))))) | (i_2_6_110_0 & i_2_6_124_0 & i_2_6_142_0))) | (i_2_6_142_0 & ((i_2_6_63_0 & ~i_2_6_84_0) | (~i_2_6_40_0 & i_2_6_110_0 & i_2_6_111_0))))) | (~i_2_6_84_0 & ((i_2_6_110_0 & ((i_2_6_34_0 & (i_2_6_111_0 | (i_2_6_32_0 & (~i_2_6_124_0 | (~i_2_6_40_0 & i_2_6_142_0))))) | (i_2_6_63_0 & i_2_6_111_0 & (i_2_6_142_0 | (~i_2_6_40_0 & ~i_2_6_124_0))))) | (i_2_6_34_0 & ((i_2_6_32_0 & ((~i_2_6_40_0 & i_2_6_111_0) | (i_2_6_63_0 & i_2_6_142_0))) | (~i_2_6_40_0 & i_2_6_63_0 & i_2_6_142_0))) | (~i_2_6_40_0 & i_2_6_63_0 & i_2_6_111_0 & i_2_6_142_0))) | (i_2_6_34_0 & ((i_2_6_63_0 & ((~i_2_6_40_0 & (i_2_6_111_0 | (i_2_6_32_0 & ~i_2_6_124_0 & (i_2_6_110_0 | i_2_6_142_0)))) | (i_2_6_110_0 & (i_2_6_111_0 | i_2_6_142_0)))) | (~i_2_6_40_0 & i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_124_0 & i_2_6_142_0))))) | (i_2_6_63_0 & ((i_2_6_34_0 & ((~i_2_6_124_0 & ((i_2_6_32_0 & ((i_2_6_62_0 & ~i_2_6_118_0) | (~i_2_6_84_0 & ~i_2_6_110_0 & ~i_2_6_142_0))) | (i_2_6_111_0 & (~i_2_6_110_0 | ~i_2_6_118_0)) | (~i_2_6_40_0 & i_2_6_62_0 & ~i_2_6_84_0 & ~i_2_6_118_0))) | (i_2_6_32_0 & ((~i_2_6_118_0 & ((i_2_6_110_0 & i_2_6_124_0) | (i_2_6_62_0 & ~i_2_6_84_0))) | (~i_2_6_84_0 & (i_2_6_111_0 | (~i_2_6_40_0 & ~i_2_6_62_0 & i_2_6_118_0 & i_2_6_124_0 & ~i_2_6_142_0))))) | (i_2_6_110_0 & ((~i_2_6_84_0 & ~i_2_6_118_0) | (~i_2_6_40_0 & i_2_6_111_0 & (~i_2_6_118_0 | (i_2_6_62_0 & ~i_2_6_84_0))))) | (i_2_6_142_0 & ((i_2_6_84_0 & i_2_6_111_0) | (i_2_6_62_0 & ~i_2_6_84_0 & ~i_2_6_118_0))))) | (~i_2_6_84_0 & ~i_2_6_118_0 & ((i_2_6_62_0 & ((~i_2_6_40_0 & i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_124_0 & i_2_6_142_0) | (i_2_6_32_0 & ((i_2_6_142_0 & (i_2_6_111_0 | (~i_2_6_40_0 & i_2_6_110_0 & ~i_2_6_124_0))) | (i_2_6_111_0 & ((i_2_6_110_0 & ~i_2_6_124_0) | (~i_2_6_40_0 & (i_2_6_110_0 | ~i_2_6_124_0)))))))) | (i_2_6_32_0 & ~i_2_6_40_0 & i_2_6_110_0 & i_2_6_111_0 & i_2_6_142_0))))) | (i_2_6_34_0 & ((i_2_6_142_0 & ((i_2_6_62_0 & ((i_2_6_40_0 & i_2_6_110_0 & i_2_6_111_0) | (i_2_6_32_0 & ~i_2_6_118_0))) | (i_2_6_32_0 & ((i_2_6_110_0 & ~i_2_6_118_0) | (~i_2_6_84_0 & ~i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_124_0))))) | (~i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_118_0 & (i_2_6_32_0 | ~i_2_6_84_0)))))) | (i_2_6_33_0 & ((~i_2_6_118_0 & ((~i_2_6_124_0 & ((~i_2_6_110_0 & ((~i_2_6_32_0 & ((~i_2_6_40_0 & i_2_6_62_0 & ~i_2_6_63_0 & ~i_2_6_84_0 & i_2_6_142_0) | (i_2_6_40_0 & i_2_6_111_0 & ~i_2_6_142_0))) | (i_2_6_32_0 & i_2_6_63_0 & ~i_2_6_84_0 & i_2_6_111_0))) | (i_2_6_62_0 & ((i_2_6_111_0 & ((~i_2_6_40_0 & (i_2_6_34_0 | (i_2_6_32_0 & i_2_6_51_0 & i_2_6_110_0 & ~i_2_6_142_0))) | (i_2_6_51_0 & i_2_6_63_0 & i_2_6_142_0))) | (~i_2_6_40_0 & ((i_2_6_142_0 & ((i_2_6_32_0 & (i_2_6_34_0 | (i_2_6_63_0 & ~i_2_6_84_0))) | (i_2_6_34_0 & i_2_6_63_0))) | (i_2_6_34_0 & ~i_2_6_84_0 & i_2_6_110_0))) | (i_2_6_32_0 & i_2_6_34_0 & (i_2_6_63_0 | i_2_6_110_0)))) | (i_2_6_34_0 & ((i_2_6_32_0 & i_2_6_142_0 & ((~i_2_6_40_0 & i_2_6_63_0) | (i_2_6_40_0 & i_2_6_110_0))) | (i_2_6_63_0 & ~i_2_6_84_0 & (~i_2_6_40_0 | i_2_6_110_0)))))) | (~i_2_6_84_0 & ((i_2_6_110_0 & ((i_2_6_32_0 & ((i_2_6_40_0 & i_2_6_124_0) | (~i_2_6_40_0 & i_2_6_62_0 & i_2_6_63_0))) | (i_2_6_34_0 & ((~i_2_6_40_0 & i_2_6_63_0) | (i_2_6_62_0 & i_2_6_142_0))) | (i_2_6_62_0 & i_2_6_111_0 & (i_2_6_142_0 | (~i_2_6_40_0 & i_2_6_63_0))) | (i_2_6_40_0 & i_2_6_63_0 & i_2_6_142_0))) | (i_2_6_34_0 & ((i_2_6_32_0 & (i_2_6_63_0 | (~i_2_6_40_0 & i_2_6_62_0))) | i_2_6_111_0 | (i_2_6_63_0 & (i_2_6_62_0 | (~i_2_6_40_0 & i_2_6_142_0))))) | (i_2_6_32_0 & ~i_2_6_40_0 & i_2_6_63_0 & ~i_2_6_110_0 & i_2_6_111_0))) | (i_2_6_34_0 & ((i_2_6_32_0 & ((i_2_6_111_0 & (i_2_6_63_0 | (~i_2_6_40_0 & i_2_6_110_0))) | (i_2_6_62_0 & ((~i_2_6_40_0 & (i_2_6_63_0 | (i_2_6_110_0 & i_2_6_142_0))) | (i_2_6_63_0 & i_2_6_110_0))))) | (i_2_6_62_0 & ((~i_2_6_40_0 & ((~i_2_6_110_0 & i_2_6_111_0) | (i_2_6_63_0 & i_2_6_110_0))) | (i_2_6_63_0 & i_2_6_110_0 & i_2_6_111_0))))))) | (i_2_6_34_0 & ((i_2_6_62_0 & ((i_2_6_110_0 & ((i_2_6_40_0 & ((i_2_6_63_0 & i_2_6_142_0) | (i_2_6_32_0 & ~i_2_6_84_0))) | (i_2_6_32_0 & (((~i_2_6_124_0 | i_2_6_142_0) & (i_2_6_63_0 | ~i_2_6_84_0)) | (i_2_6_63_0 & i_2_6_111_0))) | (~i_2_6_40_0 & i_2_6_63_0 & ~i_2_6_84_0))) | (i_2_6_32_0 & ((i_2_6_111_0 & (~i_2_6_84_0 | (~i_2_6_40_0 & i_2_6_63_0))) | (~i_2_6_40_0 & ((i_2_6_63_0 & (~i_2_6_84_0 | (~i_2_6_124_0 & i_2_6_142_0))) | (~i_2_6_84_0 & ~i_2_6_124_0 & i_2_6_142_0))) | (i_2_6_63_0 & ~i_2_6_84_0 & ~i_2_6_124_0))) | (~i_2_6_40_0 & i_2_6_63_0 & ~i_2_6_84_0 & (i_2_6_111_0 | (~i_2_6_124_0 & i_2_6_142_0))))) | (i_2_6_63_0 & ((~i_2_6_124_0 & ((i_2_6_110_0 & ((~i_2_6_40_0 & i_2_6_111_0) | (i_2_6_32_0 & ~i_2_6_84_0))) | (i_2_6_32_0 & ((~i_2_6_84_0 & i_2_6_111_0) | (~i_2_6_40_0 & i_2_6_142_0 & (~i_2_6_84_0 | i_2_6_111_0)))))) | (i_2_6_110_0 & i_2_6_111_0 & (i_2_6_142_0 | (~i_2_6_84_0 & i_2_6_124_0))))) | (~i_2_6_40_0 & ~i_2_6_84_0 & i_2_6_110_0 & i_2_6_111_0 & (~i_2_6_124_0 | i_2_6_142_0)))) | (i_2_6_62_0 & i_2_6_63_0 & i_2_6_111_0 & ((i_2_6_32_0 & ~i_2_6_40_0 & i_2_6_110_0 & ((i_2_6_124_0 & i_2_6_142_0) | (~i_2_6_84_0 & ~i_2_6_124_0))) | (~i_2_6_84_0 & i_2_6_142_0 & (~i_2_6_110_0 | ~i_2_6_124_0)))))) | (i_2_6_63_0 & ((i_2_6_34_0 & ((i_2_6_32_0 & ((i_2_6_142_0 & ((i_2_6_40_0 & ((i_2_6_62_0 & ~i_2_6_84_0) | (~i_2_6_118_0 & i_2_6_124_0))) | (i_2_6_110_0 & ((~i_2_6_84_0 & ~i_2_6_111_0) | (i_2_6_51_0 & i_2_6_62_0 & ~i_2_6_124_0))))) | (~i_2_6_84_0 & ((~i_2_6_40_0 & ((i_2_6_110_0 & i_2_6_111_0) | (i_2_6_62_0 & ~i_2_6_118_0 & ~i_2_6_124_0))) | (~i_2_6_118_0 & ((i_2_6_62_0 & i_2_6_111_0) | (i_2_6_110_0 & ~i_2_6_111_0))))) | (i_2_6_111_0 & ((i_2_6_62_0 & ~i_2_6_124_0) | (~i_2_6_118_0 & (~i_2_6_124_0 | (~i_2_6_40_0 & i_2_6_110_0))))))) | (~i_2_6_118_0 & ((i_2_6_62_0 & ((~i_2_6_40_0 & ((i_2_6_110_0 & ((i_2_6_111_0 & ~i_2_6_124_0 & i_2_6_142_0) | (~i_2_6_84_0 & (i_2_6_111_0 | (~i_2_6_124_0 & i_2_6_142_0))))) | (~i_2_6_84_0 & i_2_6_111_0 & ~i_2_6_124_0))) | (~i_2_6_84_0 & i_2_6_111_0 & (i_2_6_142_0 | (i_2_6_110_0 & ~i_2_6_124_0))))) | (i_2_6_111_0 & ~i_2_6_124_0 & i_2_6_142_0 & ~i_2_6_40_0 & ~i_2_6_84_0 & i_2_6_110_0))))) | (i_2_6_32_0 & ~i_2_6_40_0 & i_2_6_51_0 & i_2_6_62_0 & ~i_2_6_118_0 & ~i_2_6_124_0 & i_2_6_142_0 & i_2_6_110_0 & i_2_6_111_0))))) | (i_2_6_62_0 & ((~i_2_6_84_0 & ((i_2_6_34_0 & ((i_2_6_32_0 & ((~i_2_6_118_0 & ((~i_2_6_124_0 & ((~i_2_6_5_0 & ((i_2_6_40_0 & i_2_6_110_0) | (~i_2_6_63_0 & ~i_2_6_110_0 & i_2_6_142_0))) | (i_2_6_33_0 & (i_2_6_63_0 | i_2_6_110_0)) | (~i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_40_0 & i_2_6_51_0))) | (~i_2_6_40_0 & i_2_6_63_0 & (i_2_6_33_0 | (i_2_6_110_0 & i_2_6_111_0))) | (i_2_6_33_0 & (~i_2_6_51_0 | i_2_6_111_0 | (i_2_6_40_0 & i_2_6_142_0))))) | (i_2_6_63_0 & ((i_2_6_33_0 & ((~i_2_6_40_0 & (i_2_6_111_0 | (~i_2_6_124_0 & i_2_6_142_0))) | (i_2_6_110_0 & (i_2_6_111_0 | ~i_2_6_124_0)) | ~i_2_6_51_0 | (i_2_6_111_0 & ~i_2_6_124_0))) | (i_2_6_110_0 & ((~i_2_6_40_0 & ~i_2_6_51_0) | (~i_2_6_111_0 & i_2_6_142_0))) | (~i_2_6_51_0 & ~i_2_6_111_0 & (~i_2_6_124_0 | (i_2_6_118_0 & i_2_6_142_0))) | (i_2_6_51_0 & ~i_2_6_110_0 & i_2_6_111_0 & i_2_6_124_0 & i_2_6_142_0))) | (i_2_6_33_0 & ((~i_2_6_40_0 & i_2_6_111_0 & ((i_2_6_110_0 & i_2_6_142_0) | (~i_2_6_51_0 & (i_2_6_110_0 | i_2_6_142_0)))) | (~i_2_6_51_0 & i_2_6_110_0 & i_2_6_142_0))))) | (i_2_6_111_0 & ((~i_2_6_124_0 & ((i_2_6_40_0 & ((~i_2_6_51_0 & i_2_6_63_0 & i_2_6_110_0) | (i_2_6_33_0 & ~i_2_6_110_0 & ~i_2_6_118_0 & ~i_2_6_142_0))) | (i_2_6_110_0 & ((~i_2_6_40_0 & ((i_2_6_33_0 & (i_2_6_63_0 | ~i_2_6_118_0)) | (i_2_6_63_0 & ~i_2_6_118_0 & i_2_6_142_0))) | (i_2_6_33_0 & i_2_6_63_0 & i_2_6_142_0))) | (~i_2_6_32_0 & ~i_2_6_40_0 & ~i_2_6_51_0 & ~i_2_6_110_0 & ~i_2_6_118_0 & ~i_2_6_142_0))) | (i_2_6_63_0 & ((~i_2_6_118_0 & ((~i_2_6_40_0 & (i_2_6_33_0 | (~i_2_6_51_0 & i_2_6_110_0))) | (i_2_6_33_0 & (i_2_6_110_0 | i_2_6_142_0)) | (~i_2_6_51_0 & i_2_6_142_0))) | (i_2_6_33_0 & ~i_2_6_40_0 & ~i_2_6_51_0))) | (~i_2_6_118_0 & i_2_6_142_0 & i_2_6_33_0 & i_2_6_110_0))) | (i_2_6_33_0 & ((i_2_6_63_0 & ~i_2_6_118_0 & ((~i_2_6_40_0 & (i_2_6_110_0 | i_2_6_142_0)) | (i_2_6_110_0 & (~i_2_6_124_0 | i_2_6_142_0)))) | (i_2_6_40_0 & ~i_2_6_51_0 & ~i_2_6_124_0))))) | (i_2_6_33_0 & ((i_2_6_111_0 & ((~i_2_6_124_0 & ((~i_2_6_40_0 & ((i_2_6_63_0 & i_2_6_110_0 & i_2_6_32_0 & ~i_2_6_51_0) | (~i_2_6_32_0 & ~i_2_6_110_0 & i_2_6_142_0))) | (i_2_6_32_0 & ~i_2_6_118_0 & ((i_2_6_63_0 & i_2_6_142_0) | (~i_2_6_51_0 & (i_2_6_63_0 | (i_2_6_110_0 & i_2_6_142_0))))) | (~i_2_6_110_0 & i_2_6_142_0 & ~i_2_6_51_0 & i_2_6_63_0))) | (i_2_6_32_0 & ~i_2_6_51_0 & i_2_6_63_0 & ~i_2_6_118_0 & (~i_2_6_40_0 | i_2_6_110_0)))) | (~i_2_6_51_0 & i_2_6_63_0 & i_2_6_142_0 & ((i_2_6_32_0 & ~i_2_6_124_0 & (i_2_6_110_0 | ~i_2_6_118_0)) | (~i_2_6_40_0 & i_2_6_110_0 & i_2_6_124_0))))))) | (i_2_6_34_0 & ((~i_2_6_118_0 & ((i_2_6_32_0 & ((~i_2_6_124_0 & ((i_2_6_110_0 & ((i_2_6_40_0 & i_2_6_63_0 & i_2_6_142_0) | (i_2_6_33_0 & ((~i_2_6_40_0 & i_2_6_63_0) | (i_2_6_40_0 & ~i_2_6_51_0 & ~i_2_6_142_0))))) | (i_2_6_63_0 & ((~i_2_6_40_0 & i_2_6_142_0 & (i_2_6_33_0 | (~i_2_6_51_0 & i_2_6_111_0))) | (i_2_6_33_0 & (~i_2_6_51_0 | i_2_6_111_0)))) | (~i_2_6_51_0 & i_2_6_111_0 & i_2_6_33_0 & ~i_2_6_40_0))) | (~i_2_6_40_0 & ((i_2_6_33_0 & ((~i_2_6_51_0 & (i_2_6_63_0 | (i_2_6_111_0 & i_2_6_142_0))) | (i_2_6_111_0 & (i_2_6_63_0 | (i_2_6_110_0 & i_2_6_142_0))))) | (~i_2_6_51_0 & i_2_6_110_0 & ((i_2_6_63_0 & i_2_6_111_0) | (~i_2_6_63_0 & ~i_2_6_111_0 & i_2_6_142_0))))) | (i_2_6_33_0 & i_2_6_63_0 & i_2_6_142_0 & (~i_2_6_51_0 | i_2_6_111_0)))) | (i_2_6_63_0 & ((i_2_6_33_0 & ((~i_2_6_51_0 & (i_2_6_111_0 | (~i_2_6_40_0 & ~i_2_6_124_0 & i_2_6_142_0))) | (i_2_6_111_0 & ~i_2_6_124_0 & ((i_2_6_110_0 & i_2_6_142_0) | (~i_2_6_40_0 & (i_2_6_110_0 | i_2_6_142_0)))))) | (~i_2_6_40_0 & ~i_2_6_51_0 & i_2_6_110_0 & ~i_2_6_111_0 & ~i_2_6_124_0 & i_2_6_142_0))) | (i_2_6_110_0 & i_2_6_111_0 & i_2_6_142_0 & i_2_6_33_0 & ~i_2_6_51_0))) | (i_2_6_33_0 & ((~i_2_6_51_0 & ((~i_2_6_40_0 & i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_124_0 & i_2_6_142_0) | (i_2_6_63_0 & ((i_2_6_32_0 & ((~i_2_6_40_0 & (i_2_6_111_0 | (i_2_6_110_0 & ~i_2_6_124_0))) | (i_2_6_111_0 & (~i_2_6_124_0 | i_2_6_142_0)) | (~i_2_6_124_0 & i_2_6_142_0) | (i_2_6_40_0 & i_2_6_110_0 & i_2_6_124_0))) | (~i_2_6_40_0 & i_2_6_110_0 & i_2_6_142_0))))) | (i_2_6_32_0 & i_2_6_63_0 & i_2_6_111_0 & ~i_2_6_124_0 & (i_2_6_142_0 | (~i_2_6_40_0 & i_2_6_110_0))))))) | (i_2_6_33_0 & i_2_6_63_0 & i_2_6_111_0 & ~i_2_6_118_0 & i_2_6_142_0 & ((i_2_6_32_0 & ~i_2_6_51_0 & ~i_2_6_124_0 & (~i_2_6_40_0 | i_2_6_110_0)) | (i_2_6_110_0 & i_2_6_124_0 & ~i_2_6_5_0 & ~i_2_6_40_0))))) | (i_2_6_33_0 & ((i_2_6_63_0 & ((~i_2_6_51_0 & ((i_2_6_142_0 & ((~i_2_6_124_0 & ((i_2_6_32_0 & i_2_6_34_0 & ((i_2_6_110_0 & i_2_6_111_0) | (~i_2_6_40_0 & ~i_2_6_84_0))) | (~i_2_6_118_0 & ((~i_2_6_84_0 & i_2_6_111_0) | (i_2_6_40_0 & i_2_6_110_0 & ~i_2_6_111_0))))) | (i_2_6_34_0 & i_2_6_40_0 & ~i_2_6_84_0 & ~i_2_6_110_0 & i_2_6_124_0))) | (i_2_6_34_0 & ((i_2_6_111_0 & ((i_2_6_32_0 & (~i_2_6_84_0 | ~i_2_6_118_0)) | (~i_2_6_40_0 & ~i_2_6_124_0 & (~i_2_6_84_0 | i_2_6_110_0)) | (~i_2_6_84_0 & i_2_6_110_0 & i_2_6_124_0))) | (~i_2_6_40_0 & ~i_2_6_118_0 & (~i_2_6_84_0 | (i_2_6_110_0 & ~i_2_6_124_0))))) | (i_2_6_110_0 & ~i_2_6_118_0 & ~i_2_6_124_0 & ((i_2_6_32_0 & ((~i_2_6_84_0 & ~i_2_6_111_0) | (~i_2_6_40_0 & i_2_6_111_0 & ~i_2_6_142_0))) | (~i_2_6_40_0 & ~i_2_6_84_0 & i_2_6_111_0))))) | (i_2_6_34_0 & ((i_2_6_32_0 & ((i_2_6_142_0 & ((~i_2_6_40_0 & (i_2_6_111_0 | ~i_2_6_118_0) & ((~i_2_6_84_0 & ~i_2_6_124_0) | (i_2_6_110_0 & i_2_6_124_0))) | (i_2_6_111_0 & ~i_2_6_124_0 & (~i_2_6_118_0 | (~i_2_6_84_0 & i_2_6_110_0))))) | (i_2_6_110_0 & ((~i_2_6_84_0 & (~i_2_6_118_0 | (~i_2_6_40_0 & i_2_6_111_0))) | (i_2_6_111_0 & ~i_2_6_118_0))))) | (~i_2_6_84_0 & i_2_6_111_0 & ~i_2_6_118_0 & ~i_2_6_124_0 & ((i_2_6_110_0 & i_2_6_142_0) | (~i_2_6_40_0 & (i_2_6_110_0 | i_2_6_142_0)))))) | (~i_2_6_84_0 & i_2_6_110_0 & i_2_6_32_0 & ~i_2_6_40_0 & i_2_6_111_0 & ~i_2_6_118_0 & ~i_2_6_124_0 & ~i_2_6_142_0))) | (i_2_6_34_0 & i_2_6_111_0 & ((~i_2_6_84_0 & ((i_2_6_110_0 & ((i_2_6_32_0 & ~i_2_6_118_0 & (~i_2_6_40_0 | (~i_2_6_124_0 & i_2_6_142_0))) | (~i_2_6_124_0 & i_2_6_142_0 & ~i_2_6_40_0 & ~i_2_6_51_0))) | (i_2_6_32_0 & ~i_2_6_51_0 & ~i_2_6_118_0))) | (~i_2_6_118_0 & ~i_2_6_124_0 & i_2_6_142_0 & ~i_2_6_40_0 & ~i_2_6_51_0 & i_2_6_110_0))))) | (i_2_6_34_0 & ~i_2_6_51_0 & ((i_2_6_110_0 & ((~i_2_6_118_0 & ((i_2_6_32_0 & (~i_2_6_84_0 | (i_2_6_124_0 & ~i_2_6_142_0 & ~i_2_6_40_0 & i_2_6_111_0))) | (~i_2_6_84_0 & i_2_6_142_0 & ~i_2_6_40_0 & i_2_6_63_0))) | (i_2_6_118_0 & ~i_2_6_124_0 & i_2_6_142_0 & i_2_6_63_0 & ~i_2_6_84_0 & ~i_2_6_111_0))) | (i_2_6_32_0 & i_2_6_63_0 & ~i_2_6_84_0 & i_2_6_111_0 & ~i_2_6_118_0))))) | (i_2_6_34_0 & ((i_2_6_62_0 & ((~i_2_6_84_0 & ((i_2_6_32_0 & ((~i_2_6_124_0 & ((i_2_6_142_0 & ((~i_2_6_5_0 & ~i_2_6_110_0 & ((~i_2_6_33_0 & ~i_2_6_51_0) | (i_2_6_63_0 & ~i_2_6_111_0 & ~i_2_6_118_0 & i_2_6_120_0))) | (i_2_6_110_0 & ((i_2_6_33_0 & ((i_2_6_63_0 & (~i_2_6_51_0 | i_2_6_111_0)) | ~i_2_6_118_0 | (i_2_6_5_0 & i_2_6_40_0))) | (~i_2_6_40_0 & i_2_6_63_0 & i_2_6_120_0))))) | (i_2_6_111_0 & ((~i_2_6_110_0 & (i_2_6_5_0 | (~i_2_6_40_0 & ~i_2_6_51_0 & i_2_6_120_0 & ~i_2_6_142_0))) | (i_2_6_5_0 & (~i_2_6_51_0 | (i_2_6_63_0 & ~i_2_6_118_0))) | (i_2_6_33_0 & ((~i_2_6_51_0 & i_2_6_63_0) | (~i_2_6_40_0 & ((i_2_6_63_0 & i_2_6_110_0) | (~i_2_6_51_0 & ~i_2_6_142_0))))))) | (i_2_6_63_0 & ((i_2_6_33_0 & ((~i_2_6_118_0 & (~i_2_6_40_0 | i_2_6_110_0)) | (i_2_6_5_0 & (~i_2_6_51_0 | i_2_6_110_0)))) | (~i_2_6_51_0 & i_2_6_110_0 & ~i_2_6_118_0))))) | (i_2_6_110_0 & ((i_2_6_5_0 & ((~i_2_6_40_0 & ((i_2_6_111_0 & i_2_6_142_0) | (i_2_6_33_0 & i_2_6_63_0))) | (i_2_6_63_0 & ((i_2_6_124_0 & i_2_6_142_0) | (i_2_6_33_0 & (~i_2_6_51_0 | i_2_6_111_0)))))) | (i_2_6_33_0 & ((i_2_6_142_0 & ((i_2_6_63_0 & ~i_2_6_118_0) | (~i_2_6_40_0 & (~i_2_6_118_0 | (~i_2_6_51_0 & i_2_6_111_0))))) | (~i_2_6_51_0 & (~i_2_6_118_0 | (i_2_6_63_0 & i_2_6_111_0))))) | (~i_2_6_51_0 & i_2_6_63_0 & i_2_6_111_0 & ~i_2_6_118_0 & i_2_6_142_0))) | (i_2_6_33_0 & ((i_2_6_63_0 & (((i_2_6_5_0 | i_2_6_111_0) & (~i_2_6_118_0 | (~i_2_6_51_0 & (~i_2_6_40_0 | i_2_6_142_0)))) | (i_2_6_5_0 & ~i_2_6_40_0 & i_2_6_142_0))) | (i_2_6_5_0 & ~i_2_6_51_0 & i_2_6_111_0))))) | (i_2_6_33_0 & ((i_2_6_63_0 & (((~i_2_6_51_0 | (i_2_6_110_0 & ~i_2_6_124_0)) & ((i_2_6_5_0 & ~i_2_6_118_0) | (~i_2_6_40_0 & i_2_6_120_0 & i_2_6_142_0))) | (((i_2_6_111_0 & i_2_6_142_0) | (i_2_6_5_0 & i_2_6_110_0)) & ((~i_2_6_51_0 & ~i_2_6_124_0) | (~i_2_6_40_0 & ~i_2_6_118_0))) | ((~i_2_6_40_0 | i_2_6_142_0) & ((i_2_6_5_0 & ((~i_2_6_118_0 & ~i_2_6_124_0) | (~i_2_6_51_0 & i_2_6_110_0))) | (i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_118_0))) | (i_2_6_110_0 & ((i_2_6_111_0 & ((i_2_6_5_0 & (~i_2_6_40_0 | ~i_2_6_124_0)) | (~i_2_6_118_0 & ~i_2_6_124_0) | (~i_2_6_40_0 & i_2_6_142_0))) | (i_2_6_5_0 & ~i_2_6_118_0 & i_2_6_142_0))) | (~i_2_6_118_0 & ~i_2_6_124_0 & ~i_2_6_40_0 & i_2_6_111_0))) | (~i_2_6_118_0 & ((i_2_6_111_0 & (i_2_6_5_0 | (~i_2_6_51_0 & i_2_6_124_0))) | (~i_2_6_51_0 & i_2_6_142_0 & (i_2_6_110_0 | (~i_2_6_40_0 & ~i_2_6_124_0))))) | (i_2_6_5_0 & ~i_2_6_40_0 & ~i_2_6_51_0 & ((~i_2_6_124_0 & i_2_6_142_0) | (i_2_6_110_0 & (~i_2_6_124_0 | i_2_6_142_0)))))) | (i_2_6_5_0 & i_2_6_111_0 & i_2_6_142_0 & ((~i_2_6_51_0 & ~i_2_6_118_0) | (~i_2_6_40_0 & i_2_6_63_0 & i_2_6_110_0 & ~i_2_6_124_0))))) | (i_2_6_33_0 & ((i_2_6_142_0 & ((~i_2_6_124_0 & ((i_2_6_40_0 & ((i_2_6_63_0 & i_2_6_110_0 & i_2_6_5_0 & i_2_6_32_0) | (~i_2_6_51_0 & i_2_6_111_0 & ~i_2_6_118_0))) | (i_2_6_63_0 & ((~i_2_6_40_0 & ((i_2_6_5_0 & (~i_2_6_51_0 | (i_2_6_110_0 & ~i_2_6_118_0))) | (i_2_6_111_0 & (~i_2_6_51_0 | (i_2_6_32_0 & ~i_2_6_118_0))))) | (i_2_6_32_0 & i_2_6_110_0 & ((i_2_6_111_0 & ~i_2_6_118_0) | (~i_2_6_51_0 & (i_2_6_111_0 | ~i_2_6_118_0)))))))) | (~i_2_6_40_0 & ((i_2_6_5_0 & ((i_2_6_32_0 & ((i_2_6_63_0 & ~i_2_6_118_0) | (~i_2_6_51_0 & i_2_6_110_0 & i_2_6_111_0))) | (i_2_6_63_0 & ((i_2_6_110_0 & i_2_6_111_0) | (~i_2_6_51_0 & (i_2_6_110_0 | ~i_2_6_118_0)))))) | (~i_2_6_51_0 & i_2_6_110_0 & i_2_6_111_0 & (~i_2_6_118_0 | (i_2_6_32_0 & i_2_6_63_0))))) | (~i_2_6_118_0 & ((i_2_6_111_0 & ((i_2_6_5_0 & (i_2_6_32_0 | i_2_6_110_0)) | (i_2_6_32_0 & ~i_2_6_51_0 & i_2_6_63_0))) | (i_2_6_63_0 & i_2_6_110_0 & i_2_6_5_0 & ~i_2_6_51_0))))) | (i_2_6_111_0 & ((i_2_6_5_0 & ((i_2_6_32_0 & ((~i_2_6_51_0 & i_2_6_63_0 & i_2_6_110_0) | (~i_2_6_40_0 & ((~i_2_6_51_0 & i_2_6_63_0) | (~i_2_6_110_0 & ~i_2_6_118_0))))) | (~i_2_6_124_0 & ((~i_2_6_51_0 & ~i_2_6_110_0) | (i_2_6_63_0 & i_2_6_110_0 & ~i_2_6_118_0))))) | (i_2_6_32_0 & ((~i_2_6_51_0 & i_2_6_63_0 & ((~i_2_6_40_0 & (~i_2_6_118_0 | (i_2_6_110_0 & ~i_2_6_124_0))) | (~i_2_6_118_0 & (i_2_6_110_0 | ~i_2_6_124_0)))) | (~i_2_6_40_0 & i_2_6_110_0 & ~i_2_6_118_0 & i_2_6_120_0 & ~i_2_6_124_0 & ~i_2_6_142_0))) | (~i_2_6_40_0 & ~i_2_6_51_0 & i_2_6_110_0 & ~i_2_6_118_0 & ~i_2_6_124_0))) | (i_2_6_5_0 & ~i_2_6_40_0 & i_2_6_63_0 & ((i_2_6_32_0 & ~i_2_6_118_0 & (~i_2_6_51_0 | ~i_2_6_124_0)) | (~i_2_6_51_0 & i_2_6_110_0 & ~i_2_6_124_0))))) | (i_2_6_5_0 & i_2_6_32_0 & ((~i_2_6_40_0 & ((i_2_6_142_0 & ((~i_2_6_51_0 & ~i_2_6_118_0 & (i_2_6_110_0 | (~i_2_6_63_0 & ~i_2_6_124_0))) | (i_2_6_111_0 & i_2_6_118_0 & ~i_2_6_124_0))) | (i_2_6_63_0 & i_2_6_110_0 & i_2_6_111_0 & i_2_6_118_0 & ~i_2_6_124_0))) | (~i_2_6_118_0 & ((~i_2_6_51_0 & ((i_2_6_40_0 & i_2_6_63_0 & i_2_6_142_0) | (i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_124_0))) | (i_2_6_63_0 & i_2_6_110_0 & ~i_2_6_111_0 & i_2_6_120_0 & i_2_6_124_0 & i_2_6_142_0))) | (i_2_6_111_0 & i_2_6_142_0 & ~i_2_6_51_0 & i_2_6_63_0))) | (i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_40_0 & ~i_2_6_51_0 & ~i_2_6_124_0 & i_2_6_142_0 & ~i_2_6_118_0 & i_2_6_120_0))) | (~i_2_6_118_0 & ((~i_2_6_51_0 & ((~i_2_6_84_0 & ((~i_2_6_40_0 & ((~i_2_6_5_0 & ~i_2_6_63_0 & ((i_2_6_32_0 & ~i_2_6_111_0 & ~i_2_6_124_0) | (i_2_6_110_0 & i_2_6_120_0 & i_2_6_142_0))) | (i_2_6_32_0 & ((i_2_6_63_0 & i_2_6_110_0) | (i_2_6_5_0 & i_2_6_120_0 & ~i_2_6_124_0))) | (i_2_6_63_0 & ((i_2_6_33_0 & ~i_2_6_124_0) | (i_2_6_5_0 & i_2_6_110_0 & i_2_6_142_0))) | (i_2_6_5_0 & (i_2_6_33_0 | (i_2_6_111_0 & (~i_2_6_124_0 | (i_2_6_110_0 & i_2_6_120_0))))) | (i_2_6_33_0 & i_2_6_110_0 & (~i_2_6_111_0 | ~i_2_6_124_0)))) | (i_2_6_63_0 & ((i_2_6_5_0 & ((i_2_6_33_0 & i_2_6_142_0) | (i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_124_0 & ~i_2_6_142_0))) | (i_2_6_33_0 & (i_2_6_32_0 | (~i_2_6_124_0 & (i_2_6_111_0 | (i_2_6_110_0 & ~i_2_6_142_0))))))) | (i_2_6_32_0 & ((i_2_6_5_0 & (i_2_6_111_0 | i_2_6_142_0)) | (~i_2_6_124_0 & i_2_6_142_0 & i_2_6_33_0 & i_2_6_111_0))))) | (i_2_6_33_0 & ((i_2_6_63_0 & ((i_2_6_111_0 & (i_2_6_5_0 | (i_2_6_110_0 & ~i_2_6_124_0 & i_2_6_142_0))) | (~i_2_6_40_0 & ((i_2_6_32_0 & ~i_2_6_124_0 & (i_2_6_110_0 | i_2_6_142_0)) | (i_2_6_110_0 & (i_2_6_5_0 | i_2_6_142_0)))) | (i_2_6_5_0 & ((i_2_6_110_0 & ~i_2_6_124_0) | (i_2_6_32_0 & ~i_2_6_142_0 & (i_2_6_110_0 | ~i_2_6_124_0)))))) | (i_2_6_5_0 & i_2_6_32_0 & ~i_2_6_40_0 & i_2_6_110_0 & (i_2_6_111_0 | ~i_2_6_124_0)))) | (i_2_6_5_0 & i_2_6_32_0 & i_2_6_111_0 & ((~i_2_6_124_0 & i_2_6_142_0) | (~i_2_6_40_0 & i_2_6_63_0 & i_2_6_110_0))))) | (i_2_6_32_0 & ((i_2_6_5_0 & ((i_2_6_33_0 & ((i_2_6_111_0 & ((i_2_6_63_0 & ~i_2_6_124_0) | (i_2_6_124_0 & ~i_2_6_142_0 & i_2_6_40_0 & i_2_6_110_0))) | (~i_2_6_84_0 & ((i_2_6_63_0 & (~i_2_6_40_0 | (~i_2_6_124_0 & i_2_6_142_0))) | (~i_2_6_40_0 & ~i_2_6_124_0 & (i_2_6_110_0 | i_2_6_142_0)))) | (i_2_6_63_0 & i_2_6_110_0 & (~i_2_6_124_0 | (~i_2_6_40_0 & i_2_6_120_0))))) | (~i_2_6_40_0 & i_2_6_111_0 & ((~i_2_6_84_0 & i_2_6_110_0) | (~i_2_6_124_0 & ~i_2_6_142_0 & i_2_6_63_0 & ~i_2_6_110_0))))) | (i_2_6_33_0 & ((i_2_6_63_0 & ((~i_2_6_40_0 & i_2_6_110_0 & (~i_2_6_84_0 | (i_2_6_111_0 & i_2_6_142_0))) | (~i_2_6_84_0 & i_2_6_111_0 & (~i_2_6_110_0 | i_2_6_142_0)))) | (i_2_6_111_0 & ~i_2_6_124_0 & i_2_6_142_0 & ~i_2_6_40_0 & ~i_2_6_84_0 & ~i_2_6_110_0))))) | (i_2_6_33_0 & i_2_6_111_0 & ((i_2_6_142_0 & ((i_2_6_5_0 & ((~i_2_6_84_0 & ~i_2_6_124_0) | (~i_2_6_40_0 & i_2_6_63_0))) | (~i_2_6_84_0 & i_2_6_110_0 & ~i_2_6_40_0 & i_2_6_63_0))) | (i_2_6_63_0 & i_2_6_110_0 & i_2_6_5_0 & ~i_2_6_40_0))))) | (~i_2_6_84_0 & ((i_2_6_33_0 & ((i_2_6_63_0 & ((i_2_6_5_0 & ((i_2_6_32_0 & ((i_2_6_111_0 & ((i_2_6_110_0 & ~i_2_6_124_0 & i_2_6_142_0) | (~i_2_6_40_0 & ~i_2_6_110_0 & i_2_6_124_0))) | (~i_2_6_51_0 & ((i_2_6_110_0 & ~i_2_6_124_0 & i_2_6_142_0) | (~i_2_6_40_0 & (i_2_6_110_0 | (~i_2_6_124_0 & i_2_6_142_0))))))) | (i_2_6_111_0 & (~i_2_6_51_0 | (~i_2_6_40_0 & ~i_2_6_124_0 & (i_2_6_110_0 | i_2_6_142_0)))))) | (~i_2_6_51_0 & ~i_2_6_124_0 & ((~i_2_6_40_0 & ((i_2_6_111_0 & i_2_6_142_0) | (i_2_6_110_0 & ~i_2_6_142_0))) | (i_2_6_111_0 & i_2_6_142_0 & i_2_6_32_0 & i_2_6_110_0))))) | (i_2_6_5_0 & ~i_2_6_51_0 & i_2_6_110_0 & i_2_6_111_0 & i_2_6_142_0 & (~i_2_6_40_0 | (i_2_6_32_0 & ~i_2_6_124_0))))) | (i_2_6_5_0 & i_2_6_32_0 & ~i_2_6_40_0 & ~i_2_6_51_0 & i_2_6_111_0 & (i_2_6_63_0 | (i_2_6_110_0 & ~i_2_6_124_0))))) | (i_2_6_5_0 & i_2_6_33_0 & ~i_2_6_51_0 & i_2_6_63_0 & i_2_6_111_0 & ~i_2_6_124_0 & (~i_2_6_40_0 | (i_2_6_110_0 & i_2_6_142_0))))) | (i_2_6_33_0 & ((i_2_6_5_0 & ((~i_2_6_84_0 & ((~i_2_6_51_0 & ((i_2_6_62_0 & ((i_2_6_63_0 & ((~i_2_6_124_0 & ((~i_2_6_40_0 & ((i_2_6_110_0 & i_2_6_111_0) | (~i_2_6_110_0 & i_2_6_142_0))) | (i_2_6_111_0 & (~i_2_6_118_0 | i_2_6_142_0)))) | (i_2_6_110_0 & ~i_2_6_118_0 & (i_2_6_142_0 | (i_2_6_32_0 & i_2_6_111_0))))) | (~i_2_6_118_0 & i_2_6_142_0 & ~i_2_6_110_0 & i_2_6_111_0))) | (~i_2_6_118_0 & ((i_2_6_63_0 & ((i_2_6_32_0 & ((~i_2_6_40_0 & i_2_6_111_0) | (i_2_6_110_0 & ~i_2_6_111_0 & ~i_2_6_124_0))) | (i_2_6_110_0 & ((~i_2_6_124_0 & i_2_6_142_0) | (~i_2_6_40_0 & i_2_6_124_0))))) | (~i_2_6_40_0 & i_2_6_111_0 & ~i_2_6_124_0 & ~i_2_6_142_0))))) | (i_2_6_63_0 & ~i_2_6_118_0 & ((~i_2_6_40_0 & ((i_2_6_142_0 & ((i_2_6_62_0 & ((i_2_6_110_0 & ~i_2_6_124_0) | (i_2_6_120_0 & i_2_6_124_0))) | (i_2_6_110_0 & ~i_2_6_111_0 & i_2_6_120_0 & ~i_2_6_124_0))) | (i_2_6_110_0 & i_2_6_111_0 & i_2_6_32_0 & i_2_6_62_0))) | (i_2_6_32_0 & i_2_6_62_0 & i_2_6_110_0 & i_2_6_111_0 & (~i_2_6_124_0 | i_2_6_142_0)))))) | (~i_2_6_51_0 & ~i_2_6_118_0 & ((i_2_6_111_0 & ((~i_2_6_40_0 & i_2_6_63_0 & ((i_2_6_120_0 & i_2_6_142_0) | (i_2_6_32_0 & i_2_6_110_0 & ~i_2_6_124_0))) | (~i_2_6_124_0 & i_2_6_142_0 & i_2_6_62_0 & i_2_6_110_0))) | (~i_2_6_111_0 & ~i_2_6_124_0 & i_2_6_142_0 & i_2_6_40_0 & ~i_2_6_63_0 & i_2_6_110_0))))) | (i_2_6_32_0 & i_2_6_63_0 & ~i_2_6_84_0 & ~i_2_6_118_0 & ((i_2_6_142_0 & ((~i_2_6_40_0 & i_2_6_124_0 & ((~i_2_6_51_0 & i_2_6_110_0) | (i_2_6_62_0 & ~i_2_6_111_0 & i_2_6_120_0))) | (i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_124_0 & ~i_2_6_51_0 & i_2_6_62_0))) | (~i_2_6_40_0 & ~i_2_6_51_0 & i_2_6_110_0 & i_2_6_111_0 & ~i_2_6_124_0 & ~i_2_6_142_0))))) | (i_2_6_5_0 & i_2_6_32_0 & ~i_2_6_40_0 & ~i_2_6_51_0 & i_2_6_62_0 & i_2_6_63_0 & ~i_2_6_84_0 & i_2_6_110_0 & i_2_6_111_0 & i_2_6_120_0 & i_2_6_142_0);
endmodule
