module kernel_2_3 ( 
    i_2_3_29_0, i_2_3_42_0, i_2_3_43_0, i_2_3_47_0, i_2_3_55_0, i_2_3_68_0,
    i_2_3_72_0, i_2_3_77_0, i_2_3_79_0, i_2_3_86_0, i_2_3_91_0, i_2_3_99_0,
    i_2_3_138_0, i_2_3_142_0, i_2_3_143_0,
    o_2_3_0_0  );
  input  i_2_3_29_0, i_2_3_42_0, i_2_3_43_0, i_2_3_47_0, i_2_3_55_0,
    i_2_3_68_0, i_2_3_72_0, i_2_3_77_0, i_2_3_79_0, i_2_3_86_0, i_2_3_91_0,
    i_2_3_99_0, i_2_3_138_0, i_2_3_142_0, i_2_3_143_0;
  output o_2_3_0_0;
  assign o_2_3_0_0 = (~i_2_3_142_0 & ((~i_2_3_143_0 & ((~i_2_3_77_0 & ((i_2_3_68_0 & ((i_2_3_99_0 & ((~i_2_3_43_0 & ((i_2_3_79_0 & ((i_2_3_42_0 & ((i_2_3_29_0 & i_2_3_86_0 & i_2_3_91_0) | (~i_2_3_47_0 & i_2_3_55_0 & ~i_2_3_72_0 & ~i_2_3_138_0))) | (~i_2_3_42_0 & i_2_3_55_0 & i_2_3_72_0 & i_2_3_91_0))) | (i_2_3_29_0 & ~i_2_3_42_0 & ~i_2_3_47_0 & ((~i_2_3_79_0 & (i_2_3_55_0 | i_2_3_86_0)) | ~i_2_3_138_0 | (i_2_3_72_0 & i_2_3_91_0))))) | (~i_2_3_42_0 & ((i_2_3_72_0 & ((i_2_3_43_0 & ((~i_2_3_47_0 & i_2_3_86_0) | (i_2_3_29_0 & ~i_2_3_138_0))) | (i_2_3_55_0 & ((i_2_3_29_0 & (~i_2_3_138_0 | (~i_2_3_47_0 & ~i_2_3_79_0))) | (~i_2_3_47_0 & ~i_2_3_138_0) | (~i_2_3_79_0 & i_2_3_86_0))) | (i_2_3_79_0 & i_2_3_86_0 & ~i_2_3_138_0))) | (i_2_3_55_0 & ((i_2_3_29_0 & ((~i_2_3_47_0 & i_2_3_86_0) | (~i_2_3_79_0 & ~i_2_3_138_0))) | (~i_2_3_79_0 & ~i_2_3_138_0 & (~i_2_3_47_0 | i_2_3_86_0)))) | (~i_2_3_138_0 & ((~i_2_3_47_0 & (i_2_3_91_0 | (~i_2_3_79_0 & i_2_3_86_0))) | (~i_2_3_79_0 & i_2_3_86_0 & i_2_3_91_0))) | (i_2_3_86_0 & i_2_3_91_0 & i_2_3_29_0 & ~i_2_3_79_0))) | (i_2_3_29_0 & ((~i_2_3_138_0 & ((~i_2_3_79_0 & i_2_3_86_0) | (i_2_3_72_0 & (i_2_3_86_0 | (~i_2_3_47_0 & i_2_3_55_0))))) | (i_2_3_55_0 & ((i_2_3_86_0 & i_2_3_91_0) | (~i_2_3_47_0 & (i_2_3_91_0 | (~i_2_3_79_0 & i_2_3_86_0))))))) | (i_2_3_91_0 & ~i_2_3_138_0 & ((~i_2_3_47_0 & ~i_2_3_72_0 & i_2_3_79_0) | (i_2_3_72_0 & i_2_3_86_0))))) | (~i_2_3_138_0 & ((i_2_3_29_0 & ((i_2_3_43_0 & ((~i_2_3_42_0 & i_2_3_72_0 & ~i_2_3_79_0) | (i_2_3_55_0 & ~i_2_3_72_0 & i_2_3_79_0 & i_2_3_86_0 & ~i_2_3_99_0))) | (~i_2_3_79_0 & (((i_2_3_55_0 | i_2_3_86_0) & ((~i_2_3_43_0 & ~i_2_3_47_0) | i_2_3_91_0 | (~i_2_3_42_0 & i_2_3_72_0))) | (~i_2_3_47_0 & ((~i_2_3_42_0 & ~i_2_3_43_0) | (i_2_3_55_0 & i_2_3_72_0))) | (i_2_3_55_0 & i_2_3_72_0 & i_2_3_86_0))) | (~i_2_3_42_0 & (((i_2_3_55_0 | i_2_3_86_0) & (~i_2_3_47_0 | i_2_3_91_0)) | (i_2_3_55_0 & i_2_3_86_0))) | (~i_2_3_47_0 & i_2_3_72_0 & i_2_3_91_0))) | (~i_2_3_47_0 & (((i_2_3_55_0 | i_2_3_86_0) & ((i_2_3_72_0 & ((~i_2_3_42_0 & ~i_2_3_79_0) | (~i_2_3_43_0 & i_2_3_91_0))) | (~i_2_3_79_0 & i_2_3_91_0))) | (i_2_3_86_0 & ((~i_2_3_42_0 & (i_2_3_55_0 | i_2_3_91_0)) | (i_2_3_55_0 & i_2_3_72_0 & ~i_2_3_79_0))) | (~i_2_3_42_0 & ~i_2_3_79_0 & i_2_3_91_0))) | (~i_2_3_42_0 & ((~i_2_3_79_0 & ((i_2_3_55_0 & (i_2_3_91_0 | (i_2_3_72_0 & i_2_3_86_0))) | (i_2_3_72_0 & i_2_3_86_0 & i_2_3_91_0))) | (i_2_3_55_0 & i_2_3_86_0 & i_2_3_91_0))) | (i_2_3_86_0 & i_2_3_91_0 & i_2_3_55_0 & ~i_2_3_79_0))) | (~i_2_3_42_0 & ((i_2_3_91_0 & ((i_2_3_29_0 & ((i_2_3_72_0 & ((~i_2_3_47_0 & i_2_3_86_0) | (~i_2_3_43_0 & i_2_3_55_0 & ~i_2_3_79_0))) | (i_2_3_86_0 & (~i_2_3_47_0 | i_2_3_55_0) & (~i_2_3_43_0 | ~i_2_3_79_0)))) | (~i_2_3_43_0 & ~i_2_3_47_0 & i_2_3_86_0 & (i_2_3_55_0 | (i_2_3_72_0 & ~i_2_3_79_0))))) | (i_2_3_29_0 & ~i_2_3_47_0 & i_2_3_55_0 & i_2_3_86_0 & (i_2_3_72_0 | ~i_2_3_79_0)))) | (i_2_3_55_0 & i_2_3_86_0 & i_2_3_91_0 & i_2_3_29_0 & ~i_2_3_47_0))) | (i_2_3_29_0 & ((i_2_3_91_0 & ((i_2_3_43_0 & ~i_2_3_68_0 & ((~i_2_3_47_0 & ~i_2_3_138_0) | (~i_2_3_42_0 & i_2_3_55_0 & ~i_2_3_79_0))) | (~i_2_3_42_0 & ((~i_2_3_47_0 & ((i_2_3_55_0 & ((i_2_3_72_0 & i_2_3_99_0) | (~i_2_3_72_0 & i_2_3_79_0 & ~i_2_3_99_0))) | (i_2_3_99_0 & (~i_2_3_138_0 | (i_2_3_72_0 & i_2_3_86_0))) | (i_2_3_72_0 & (~i_2_3_138_0 | (~i_2_3_43_0 & ~i_2_3_79_0 & ~i_2_3_99_0))))) | (i_2_3_55_0 & ((~i_2_3_79_0 & (~i_2_3_138_0 | (i_2_3_86_0 & i_2_3_99_0))) | (i_2_3_99_0 & ~i_2_3_138_0))) | (i_2_3_86_0 & ~i_2_3_138_0 & (~i_2_3_79_0 | i_2_3_99_0)))) | (~i_2_3_138_0 & ((i_2_3_72_0 & ((i_2_3_55_0 & i_2_3_86_0) | (~i_2_3_79_0 & i_2_3_99_0))) | (i_2_3_55_0 & (~i_2_3_47_0 | (i_2_3_86_0 & (~i_2_3_79_0 | i_2_3_99_0)))))) | (~i_2_3_47_0 & i_2_3_72_0 & ~i_2_3_79_0 & (i_2_3_55_0 | (i_2_3_86_0 & ~i_2_3_99_0))))) | (~i_2_3_138_0 & ((i_2_3_86_0 & ((~i_2_3_47_0 & ((~i_2_3_42_0 & (~i_2_3_79_0 | (i_2_3_43_0 & ~i_2_3_72_0))) | (i_2_3_72_0 & (i_2_3_99_0 | (i_2_3_43_0 & ~i_2_3_79_0))) | i_2_3_55_0 | (~i_2_3_43_0 & i_2_3_99_0))) | (i_2_3_55_0 & ((~i_2_3_42_0 & ((~i_2_3_79_0 & i_2_3_99_0) | ((~i_2_3_79_0 | i_2_3_99_0) & (~i_2_3_43_0 | i_2_3_72_0)))) | (i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_99_0))))) | (~i_2_3_42_0 & ((i_2_3_55_0 & ((~i_2_3_43_0 & i_2_3_72_0 & (~i_2_3_47_0 | (~i_2_3_79_0 & i_2_3_99_0))) | (~i_2_3_47_0 & (~i_2_3_79_0 | i_2_3_99_0)))) | (~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_47_0 & i_2_3_72_0))) | (~i_2_3_47_0 & i_2_3_55_0 & i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_99_0))) | (~i_2_3_42_0 & ~i_2_3_47_0 & i_2_3_55_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0))) | (i_2_3_86_0 & ((i_2_3_72_0 & ((i_2_3_99_0 & ((i_2_3_91_0 & ((~i_2_3_42_0 & (i_2_3_55_0 | (~i_2_3_29_0 & i_2_3_47_0 & ~i_2_3_68_0 & ~i_2_3_79_0))) | (i_2_3_55_0 & (~i_2_3_47_0 | (~i_2_3_79_0 & ~i_2_3_138_0))))) | (~i_2_3_43_0 & ~i_2_3_47_0 & ~i_2_3_68_0 & ~i_2_3_79_0 & ~i_2_3_138_0))) | (~i_2_3_47_0 & ((i_2_3_55_0 & ((~i_2_3_42_0 & ((i_2_3_43_0 & i_2_3_91_0) | (~i_2_3_43_0 & ~i_2_3_138_0))) | (~i_2_3_43_0 & ~i_2_3_79_0 & i_2_3_91_0))) | (~i_2_3_42_0 & i_2_3_91_0 & ~i_2_3_138_0))))) | (~i_2_3_42_0 & ((~i_2_3_138_0 & ((~i_2_3_47_0 & ((i_2_3_43_0 & (i_2_3_91_0 | (i_2_3_55_0 & ~i_2_3_72_0))) | ((i_2_3_55_0 | i_2_3_91_0) & (~i_2_3_79_0 | i_2_3_99_0)))) | (i_2_3_55_0 & i_2_3_91_0 & (~i_2_3_79_0 | i_2_3_99_0)))) | (~i_2_3_47_0 & i_2_3_55_0 & ~i_2_3_79_0 & i_2_3_91_0))))) | (~i_2_3_47_0 & ((i_2_3_55_0 & ((~i_2_3_42_0 & ((i_2_3_72_0 & ((i_2_3_91_0 & ~i_2_3_138_0) | (~i_2_3_79_0 & ((i_2_3_99_0 & ~i_2_3_138_0) | (~i_2_3_43_0 & i_2_3_91_0 & ~i_2_3_99_0))))) | (i_2_3_91_0 & i_2_3_99_0 & ~i_2_3_138_0))) | (i_2_3_91_0 & ~i_2_3_138_0 & ~i_2_3_72_0 & ~i_2_3_79_0))) | (i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_91_0 & i_2_3_99_0 & ~i_2_3_138_0))) | (~i_2_3_42_0 & i_2_3_43_0 & i_2_3_55_0 & i_2_3_72_0 & i_2_3_91_0 & ~i_2_3_138_0))) | (~i_2_3_138_0 & ((i_2_3_91_0 & ((i_2_3_68_0 & ((i_2_3_43_0 & ((~i_2_3_47_0 & ~i_2_3_86_0 & i_2_3_99_0) | (i_2_3_86_0 & ~i_2_3_99_0 & ~i_2_3_42_0 & i_2_3_72_0))) | ((i_2_3_29_0 | ~i_2_3_47_0) & ((i_2_3_86_0 & ((i_2_3_55_0 & i_2_3_72_0) | (~i_2_3_42_0 & (i_2_3_72_0 | ~i_2_3_79_0)))) | (i_2_3_55_0 & ~i_2_3_72_0 & i_2_3_99_0))) | (~i_2_3_47_0 & (((~i_2_3_42_0 | ~i_2_3_79_0) & (i_2_3_29_0 | (i_2_3_86_0 & i_2_3_99_0))) | (~i_2_3_42_0 & i_2_3_55_0 & ~i_2_3_79_0) | (i_2_3_72_0 & ((~i_2_3_42_0 & i_2_3_55_0) | (i_2_3_29_0 & (i_2_3_55_0 | i_2_3_86_0)))))) | (i_2_3_29_0 & ((i_2_3_55_0 & ~i_2_3_79_0 & i_2_3_86_0) | (~i_2_3_42_0 & i_2_3_99_0))) | (i_2_3_72_0 & ((~i_2_3_42_0 & ((i_2_3_55_0 & i_2_3_86_0) | (i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_99_0))) | (i_2_3_55_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0))) | (~i_2_3_42_0 & i_2_3_55_0 & ~i_2_3_79_0 & i_2_3_86_0))) | (~i_2_3_47_0 & ((i_2_3_29_0 & ((~i_2_3_42_0 & (i_2_3_55_0 | i_2_3_86_0)) | (~i_2_3_72_0 & (~i_2_3_79_0 | (~i_2_3_43_0 & i_2_3_55_0))) | (i_2_3_72_0 & i_2_3_99_0) | (i_2_3_77_0 & ~i_2_3_79_0))) | (i_2_3_72_0 & ((i_2_3_86_0 & (~i_2_3_79_0 | i_2_3_99_0) & (i_2_3_55_0 | (~i_2_3_42_0 & ~i_2_3_43_0))) | (~i_2_3_42_0 & i_2_3_55_0 & (~i_2_3_79_0 | (~i_2_3_43_0 & i_2_3_99_0))))) | (~i_2_3_42_0 & i_2_3_86_0 & (i_2_3_55_0 | (~i_2_3_79_0 & i_2_3_99_0))) | (i_2_3_55_0 & ~i_2_3_79_0 & i_2_3_99_0))) | (i_2_3_29_0 & ((~i_2_3_42_0 & ((~i_2_3_43_0 & ((i_2_3_55_0 & i_2_3_86_0) | (i_2_3_72_0 & i_2_3_77_0 & i_2_3_99_0))) | (~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0) | (i_2_3_55_0 & ((i_2_3_86_0 & i_2_3_99_0) | (~i_2_3_79_0 & (i_2_3_86_0 | i_2_3_99_0)))))) | (i_2_3_55_0 & ~i_2_3_79_0 & i_2_3_86_0 & (i_2_3_72_0 | i_2_3_99_0)))) | (~i_2_3_42_0 & i_2_3_55_0 & ~i_2_3_79_0 & i_2_3_99_0 & (i_2_3_72_0 | (~i_2_3_43_0 & i_2_3_86_0))))) | (~i_2_3_47_0 & ((i_2_3_68_0 & ((~i_2_3_79_0 & ((i_2_3_99_0 & ((i_2_3_72_0 & ((i_2_3_55_0 & i_2_3_86_0) | (~i_2_3_42_0 & (i_2_3_55_0 | i_2_3_86_0)))) | (i_2_3_43_0 & (~i_2_3_55_0 | i_2_3_86_0)) | (i_2_3_29_0 & i_2_3_55_0))) | (i_2_3_55_0 & ((i_2_3_29_0 & (~i_2_3_42_0 | i_2_3_86_0)) | (~i_2_3_42_0 & i_2_3_86_0))))) | (~i_2_3_42_0 & ((i_2_3_29_0 & (i_2_3_55_0 | i_2_3_86_0) & (i_2_3_72_0 | i_2_3_99_0)) | (i_2_3_55_0 & i_2_3_86_0 & (i_2_3_99_0 | (~i_2_3_43_0 & i_2_3_72_0))))) | (i_2_3_72_0 & i_2_3_86_0 & i_2_3_29_0 & i_2_3_55_0))) | (i_2_3_29_0 & ((~i_2_3_43_0 & ((i_2_3_99_0 & ((~i_2_3_42_0 & i_2_3_55_0 & i_2_3_72_0) | (~i_2_3_68_0 & ~i_2_3_79_0 & i_2_3_86_0))) | (i_2_3_55_0 & ((~i_2_3_42_0 & (i_2_3_86_0 | (i_2_3_72_0 & ~i_2_3_79_0))) | (i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_86_0))))) | (i_2_3_86_0 & ((i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_99_0) | (~i_2_3_42_0 & i_2_3_55_0 & (i_2_3_72_0 | i_2_3_99_0)))) | (~i_2_3_42_0 & i_2_3_55_0 & ~i_2_3_79_0 & i_2_3_99_0))) | (~i_2_3_42_0 & i_2_3_55_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0 & (~i_2_3_43_0 | i_2_3_72_0)))) | (i_2_3_29_0 & ((~i_2_3_42_0 & i_2_3_55_0 & ((i_2_3_86_0 & ((~i_2_3_43_0 & ((~i_2_3_79_0 & i_2_3_99_0) | (i_2_3_68_0 & i_2_3_72_0))) | (i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_99_0) | (i_2_3_68_0 & (~i_2_3_79_0 | i_2_3_99_0)))) | (~i_2_3_79_0 & i_2_3_99_0 & i_2_3_68_0 & i_2_3_72_0))) | (~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0 & i_2_3_68_0 & i_2_3_72_0))) | (~i_2_3_42_0 & ~i_2_3_43_0 & i_2_3_55_0 & i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0))) | (i_2_3_29_0 & ((i_2_3_91_0 & ((~i_2_3_42_0 & ((~i_2_3_79_0 & ((i_2_3_99_0 & ((i_2_3_43_0 & (i_2_3_72_0 | (~i_2_3_47_0 & i_2_3_86_0))) | (i_2_3_55_0 & i_2_3_68_0 & ~i_2_3_72_0))) | (i_2_3_55_0 & i_2_3_72_0 & i_2_3_86_0) | (~i_2_3_47_0 & i_2_3_68_0 & ((i_2_3_72_0 & i_2_3_86_0) | (~i_2_3_43_0 & (i_2_3_55_0 | i_2_3_86_0)))))) | (i_2_3_68_0 & ((~i_2_3_47_0 & ((i_2_3_86_0 & i_2_3_99_0) | (i_2_3_55_0 & (i_2_3_86_0 | i_2_3_99_0)))) | (i_2_3_55_0 & i_2_3_72_0 & i_2_3_86_0 & i_2_3_99_0))))) | (~i_2_3_47_0 & ((~i_2_3_79_0 & ((~i_2_3_43_0 & ((i_2_3_55_0 & i_2_3_86_0) | (i_2_3_72_0 & i_2_3_77_0 & i_2_3_99_0))) | (i_2_3_55_0 & i_2_3_72_0 & i_2_3_86_0) | (i_2_3_68_0 & ~i_2_3_72_0 & i_2_3_99_0))) | (i_2_3_55_0 & i_2_3_86_0 & i_2_3_99_0 & (i_2_3_43_0 | i_2_3_68_0 | ~i_2_3_72_0)))))) | (~i_2_3_42_0 & ~i_2_3_47_0 & i_2_3_55_0 & i_2_3_68_0 & i_2_3_86_0 & ((~i_2_3_79_0 & i_2_3_99_0) | (i_2_3_72_0 & (~i_2_3_79_0 | i_2_3_99_0)))))) | (~i_2_3_47_0 & i_2_3_55_0 & i_2_3_72_0 & i_2_3_86_0 & i_2_3_91_0 & ((~i_2_3_79_0 & i_2_3_99_0) | (~i_2_3_42_0 & i_2_3_68_0 & (~i_2_3_79_0 | i_2_3_99_0)))))) | (i_2_3_29_0 & ((~i_2_3_42_0 & ((i_2_3_72_0 & ((~i_2_3_79_0 & ((~i_2_3_55_0 & ((~i_2_3_47_0 & ~i_2_3_68_0 & ~i_2_3_86_0 & i_2_3_91_0 & ~i_2_3_99_0) | (~i_2_3_43_0 & ~i_2_3_77_0 & i_2_3_86_0 & ~i_2_3_138_0 & i_2_3_143_0))) | (i_2_3_86_0 & ((~i_2_3_138_0 & ((~i_2_3_43_0 & (i_2_3_91_0 | (i_2_3_68_0 & i_2_3_143_0))) | (i_2_3_55_0 & (~i_2_3_47_0 | (~i_2_3_77_0 & i_2_3_99_0))))) | (i_2_3_68_0 & ((~i_2_3_47_0 & ((i_2_3_55_0 & (~i_2_3_77_0 | i_2_3_99_0)) | (~i_2_3_77_0 & i_2_3_91_0))) | (i_2_3_77_0 & i_2_3_91_0 & i_2_3_99_0 & i_2_3_143_0))) | (~i_2_3_77_0 & i_2_3_91_0 & (i_2_3_55_0 | (i_2_3_43_0 & ~i_2_3_68_0 & i_2_3_138_0))))) | (~i_2_3_47_0 & ((~i_2_3_77_0 & ((~i_2_3_43_0 & ((i_2_3_68_0 & i_2_3_91_0 & i_2_3_99_0) | (i_2_3_55_0 & ~i_2_3_138_0))) | (i_2_3_55_0 & i_2_3_91_0 & i_2_3_99_0))) | (i_2_3_55_0 & i_2_3_68_0 & ~i_2_3_138_0))) | (~i_2_3_138_0 & ((i_2_3_55_0 & i_2_3_91_0) | (i_2_3_99_0 & i_2_3_143_0 & i_2_3_68_0 & ~i_2_3_77_0))))) | (~i_2_3_138_0 & ((i_2_3_68_0 & ((i_2_3_91_0 & (i_2_3_55_0 | (~i_2_3_77_0 & i_2_3_143_0))) | (i_2_3_55_0 & (~i_2_3_77_0 | i_2_3_99_0) & (~i_2_3_47_0 | (~i_2_3_43_0 & i_2_3_86_0))) | (~i_2_3_47_0 & ((~i_2_3_77_0 & i_2_3_86_0) | (i_2_3_99_0 & i_2_3_143_0 & ~i_2_3_43_0 & i_2_3_77_0))))) | (~i_2_3_47_0 & ((~i_2_3_43_0 & (i_2_3_55_0 | i_2_3_86_0) & (i_2_3_91_0 | (~i_2_3_77_0 & i_2_3_99_0))) | (i_2_3_55_0 & i_2_3_86_0 & (~i_2_3_77_0 | i_2_3_99_0)))) | (i_2_3_91_0 & ((i_2_3_55_0 & (~i_2_3_77_0 | (i_2_3_99_0 & i_2_3_143_0))) | (~i_2_3_77_0 & i_2_3_86_0 & (~i_2_3_43_0 | (i_2_3_79_0 & ~i_2_3_99_0))))))) | (~i_2_3_47_0 & ((i_2_3_55_0 & ((i_2_3_91_0 & ((~i_2_3_43_0 & ((i_2_3_86_0 & i_2_3_99_0) | (i_2_3_68_0 & ~i_2_3_77_0))) | (i_2_3_68_0 & i_2_3_86_0))) | (i_2_3_86_0 & i_2_3_99_0 & i_2_3_68_0 & ~i_2_3_77_0))) | (i_2_3_68_0 & ~i_2_3_77_0 & i_2_3_86_0 & i_2_3_91_0 & i_2_3_99_0))))) | (~i_2_3_138_0 & ((i_2_3_91_0 & ((i_2_3_43_0 & ((~i_2_3_47_0 & i_2_3_68_0 & i_2_3_77_0) | (i_2_3_55_0 & ~i_2_3_79_0 & ~i_2_3_86_0))) | (i_2_3_55_0 & ((i_2_3_86_0 & ((~i_2_3_43_0 & (~i_2_3_79_0 | i_2_3_99_0)) | (~i_2_3_79_0 & i_2_3_99_0) | i_2_3_68_0 | ~i_2_3_77_0)) | (~i_2_3_47_0 & (~i_2_3_77_0 | i_2_3_99_0)) | (i_2_3_68_0 & ~i_2_3_79_0))) | (i_2_3_68_0 & ((~i_2_3_43_0 & ((~i_2_3_47_0 & ~i_2_3_72_0) | (~i_2_3_77_0 & ~i_2_3_79_0))) | (~i_2_3_77_0 & i_2_3_86_0 & i_2_3_99_0))) | (i_2_3_86_0 & i_2_3_99_0 & (~i_2_3_47_0 | (~i_2_3_77_0 & ~i_2_3_79_0))))) | (i_2_3_55_0 & (((~i_2_3_79_0 | i_2_3_99_0) & ((~i_2_3_47_0 & ((~i_2_3_43_0 & i_2_3_86_0) | (i_2_3_68_0 & ~i_2_3_77_0))) | (i_2_3_68_0 & ~i_2_3_77_0 & i_2_3_86_0))) | (i_2_3_86_0 & ((i_2_3_68_0 & (~i_2_3_47_0 | (~i_2_3_79_0 & i_2_3_99_0))) | (i_2_3_99_0 & ((~i_2_3_47_0 & (~i_2_3_77_0 | ~i_2_3_79_0)) | (~i_2_3_43_0 & ~i_2_3_77_0 & ~i_2_3_79_0))))) | (~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_47_0 & ~i_2_3_77_0))) | (~i_2_3_47_0 & ((i_2_3_86_0 & ((i_2_3_68_0 & ((~i_2_3_72_0 & ~i_2_3_79_0) | (~i_2_3_77_0 & i_2_3_99_0))) | (~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_99_0))) | (i_2_3_68_0 & i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_99_0 & i_2_3_143_0))))) | (i_2_3_68_0 & ((i_2_3_91_0 & (((~i_2_3_79_0 | i_2_3_99_0) & ((~i_2_3_77_0 & ((~i_2_3_47_0 & i_2_3_55_0) | (~i_2_3_43_0 & i_2_3_86_0 & (~i_2_3_47_0 | i_2_3_55_0)))) | (~i_2_3_47_0 & i_2_3_55_0 & i_2_3_86_0))) | (~i_2_3_47_0 & ~i_2_3_79_0 & i_2_3_99_0 & (i_2_3_55_0 | i_2_3_86_0)))) | (~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_47_0 & i_2_3_55_0 & ~i_2_3_77_0))) | (~i_2_3_47_0 & i_2_3_55_0 & ~i_2_3_77_0 & i_2_3_86_0 & i_2_3_91_0))) | (~i_2_3_138_0 & ((i_2_3_91_0 & ((~i_2_3_47_0 & ((~i_2_3_43_0 & ((i_2_3_68_0 & ~i_2_3_72_0 & i_2_3_86_0) | (~i_2_3_79_0 & i_2_3_143_0))) | (i_2_3_55_0 & (i_2_3_86_0 | (i_2_3_68_0 & ~i_2_3_77_0))) | (~i_2_3_77_0 & i_2_3_86_0) | (~i_2_3_68_0 & ((~i_2_3_79_0 & i_2_3_86_0) | (i_2_3_72_0 & ~i_2_3_77_0 & i_2_3_79_0 & i_2_3_99_0))))) | (i_2_3_55_0 & ((~i_2_3_77_0 & ((~i_2_3_43_0 & ((~i_2_3_79_0 & i_2_3_99_0) | (i_2_3_68_0 & (i_2_3_72_0 | i_2_3_86_0)))) | (i_2_3_86_0 & i_2_3_99_0 & (i_2_3_72_0 | ~i_2_3_79_0)))) | (i_2_3_72_0 & i_2_3_99_0 & ((~i_2_3_43_0 & i_2_3_86_0) | (i_2_3_68_0 & i_2_3_79_0 & i_2_3_143_0))))) | (i_2_3_68_0 & ((i_2_3_143_0 & ((i_2_3_72_0 & ((i_2_3_86_0 & i_2_3_99_0) | (i_2_3_77_0 & ~i_2_3_79_0 & ~i_2_3_99_0))) | (~i_2_3_79_0 & ((i_2_3_86_0 & i_2_3_99_0) | (i_2_3_43_0 & i_2_3_47_0 & ~i_2_3_77_0))))) | (~i_2_3_43_0 & ~i_2_3_79_0 & i_2_3_99_0))))) | (~i_2_3_47_0 & ((i_2_3_72_0 & ((i_2_3_68_0 & ((i_2_3_55_0 & i_2_3_86_0 & (~i_2_3_77_0 | ~i_2_3_79_0)) | (~i_2_3_79_0 & i_2_3_99_0 & (~i_2_3_55_0 | ~i_2_3_77_0)))) | (i_2_3_55_0 & ~i_2_3_77_0 & i_2_3_86_0 & (~i_2_3_79_0 | i_2_3_99_0)))) | (i_2_3_55_0 & i_2_3_86_0 & ((~i_2_3_77_0 & (~i_2_3_43_0 | (~i_2_3_79_0 & i_2_3_99_0))) | (i_2_3_68_0 & i_2_3_99_0))))))) | (~i_2_3_77_0 & ((~i_2_3_79_0 & ((i_2_3_72_0 & ((i_2_3_91_0 & ((i_2_3_86_0 & ((~i_2_3_43_0 & ((~i_2_3_47_0 & i_2_3_99_0) | (i_2_3_55_0 & ~i_2_3_99_0))) | (~i_2_3_47_0 & i_2_3_68_0 & i_2_3_99_0) | (i_2_3_55_0 & ~i_2_3_68_0 & ~i_2_3_99_0))) | (~i_2_3_47_0 & i_2_3_55_0 & i_2_3_68_0 & i_2_3_99_0))) | (~i_2_3_43_0 & ~i_2_3_47_0 & i_2_3_55_0 & ~i_2_3_68_0 & i_2_3_86_0))) | (i_2_3_86_0 & i_2_3_91_0 & ~i_2_3_47_0 & i_2_3_55_0))) | (i_2_3_86_0 & i_2_3_91_0 & i_2_3_99_0 & ~i_2_3_47_0 & i_2_3_55_0 & i_2_3_68_0))) | (i_2_3_86_0 & i_2_3_91_0 & i_2_3_99_0 & ~i_2_3_47_0 & i_2_3_55_0 & ~i_2_3_79_0))) | (~i_2_3_47_0 & ((i_2_3_91_0 & ((~i_2_3_138_0 & ((i_2_3_55_0 & ((i_2_3_43_0 & ((~i_2_3_68_0 & ~i_2_3_77_0 & ~i_2_3_79_0) | (~i_2_3_42_0 & i_2_3_68_0 & ~i_2_3_99_0))) | (i_2_3_86_0 & ((~i_2_3_43_0 & ((~i_2_3_42_0 & i_2_3_99_0) | (i_2_3_68_0 & ~i_2_3_72_0))) | (i_2_3_68_0 & (~i_2_3_42_0 | ~i_2_3_79_0)) | (~i_2_3_42_0 & (~i_2_3_79_0 | (i_2_3_72_0 & i_2_3_99_0))) | ~i_2_3_77_0 | (~i_2_3_79_0 & i_2_3_99_0))) | (~i_2_3_42_0 & ((i_2_3_68_0 & (~i_2_3_77_0 | (i_2_3_72_0 & ~i_2_3_79_0))) | (i_2_3_72_0 & ~i_2_3_77_0 & i_2_3_99_0))) | (~i_2_3_43_0 & i_2_3_72_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & ~i_2_3_99_0 & i_2_3_143_0))) | (i_2_3_86_0 & ((i_2_3_72_0 & ((~i_2_3_79_0 & ((~i_2_3_43_0 & ((~i_2_3_42_0 & i_2_3_99_0) | (~i_2_3_77_0 & i_2_3_143_0))) | (~i_2_3_42_0 & (i_2_3_68_0 | ~i_2_3_77_0)))) | (~i_2_3_42_0 & i_2_3_99_0 & (i_2_3_68_0 | ~i_2_3_77_0)))) | (~i_2_3_42_0 & ~i_2_3_77_0 & ((~i_2_3_79_0 & i_2_3_99_0) | (i_2_3_68_0 & (~i_2_3_79_0 | i_2_3_99_0)))))) | (i_2_3_68_0 & ~i_2_3_79_0 & i_2_3_99_0 & ((~i_2_3_77_0 & i_2_3_143_0) | (~i_2_3_42_0 & ~i_2_3_72_0))))) | (~i_2_3_42_0 & i_2_3_68_0 & ((~i_2_3_77_0 & ((~i_2_3_43_0 & ((~i_2_3_79_0 & ((i_2_3_55_0 & (i_2_3_86_0 | (i_2_3_72_0 & i_2_3_99_0))) | (i_2_3_72_0 & i_2_3_86_0 & i_2_3_99_0))) | (i_2_3_55_0 & i_2_3_86_0 & i_2_3_99_0))) | (~i_2_3_79_0 & i_2_3_86_0 & i_2_3_55_0 & i_2_3_72_0))) | (i_2_3_55_0 & i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0))) | (i_2_3_55_0 & ~i_2_3_68_0 & i_2_3_72_0 & i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_77_0 & ~i_2_3_79_0))) | (~i_2_3_138_0 & ((i_2_3_55_0 & ((i_2_3_86_0 & ((i_2_3_68_0 & ((i_2_3_72_0 & ((~i_2_3_42_0 & (~i_2_3_77_0 | (~i_2_3_43_0 & ~i_2_3_79_0))) | (i_2_3_99_0 & i_2_3_143_0 & ~i_2_3_43_0 & i_2_3_79_0))) | (~i_2_3_42_0 & ~i_2_3_79_0 & (~i_2_3_77_0 | i_2_3_99_0)) | (~i_2_3_72_0 & ~i_2_3_77_0 & i_2_3_99_0))) | (~i_2_3_77_0 & ~i_2_3_79_0 & ((i_2_3_72_0 & i_2_3_99_0) | (~i_2_3_42_0 & (i_2_3_99_0 | (i_2_3_43_0 & ~i_2_3_72_0))))))) | (~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_42_0 & i_2_3_68_0 & i_2_3_72_0))) | (i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & ~i_2_3_42_0 & i_2_3_68_0 & i_2_3_72_0))))) | (i_2_3_55_0 & ((i_2_3_91_0 & ((i_2_3_99_0 & ((~i_2_3_138_0 & ((~i_2_3_79_0 & ((~i_2_3_42_0 & ((~i_2_3_77_0 & i_2_3_86_0) | (~i_2_3_43_0 & i_2_3_72_0 & ~i_2_3_86_0))) | (~i_2_3_43_0 & i_2_3_68_0 & ~i_2_3_77_0))) | (i_2_3_68_0 & i_2_3_79_0 & ((~i_2_3_72_0 & ~i_2_3_77_0) | (i_2_3_72_0 & i_2_3_86_0 & i_2_3_143_0))))) | (~i_2_3_42_0 & i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_77_0 & i_2_3_86_0))) | (~i_2_3_42_0 & i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_86_0 & ~i_2_3_138_0))) | (~i_2_3_42_0 & i_2_3_68_0 & i_2_3_72_0 & i_2_3_99_0 & ~i_2_3_138_0 & ~i_2_3_77_0 & i_2_3_86_0))) | (~i_2_3_42_0 & i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_77_0 & i_2_3_79_0 & i_2_3_86_0 & i_2_3_91_0 & ~i_2_3_99_0 & ~i_2_3_138_0 & i_2_3_143_0))) | (~i_2_3_47_0 & ((i_2_3_91_0 & ((~i_2_3_42_0 & ((i_2_3_55_0 & ((~i_2_3_143_0 & ((i_2_3_72_0 & ((~i_2_3_43_0 & ((i_2_3_29_0 & i_2_3_86_0 & ~i_2_3_99_0) | (~i_2_3_68_0 & ~i_2_3_77_0 & i_2_3_99_0 & i_2_3_142_0))) | (i_2_3_99_0 & ((i_2_3_86_0 & ~i_2_3_138_0) | (i_2_3_29_0 & i_2_3_68_0 & ~i_2_3_77_0))) | (~i_2_3_79_0 & ((i_2_3_29_0 & (i_2_3_43_0 | ~i_2_3_77_0)) | (~i_2_3_77_0 & (~i_2_3_138_0 | (i_2_3_86_0 & ~i_2_3_99_0))) | (~i_2_3_138_0 & (i_2_3_68_0 | i_2_3_86_0)))) | (i_2_3_68_0 & ~i_2_3_77_0 & ~i_2_3_138_0))) | (~i_2_3_77_0 & ((i_2_3_29_0 & (~i_2_3_138_0 | (i_2_3_43_0 & ~i_2_3_99_0))) | (~i_2_3_72_0 & ((i_2_3_68_0 & ~i_2_3_79_0 & i_2_3_99_0) | (i_2_3_43_0 & ~i_2_3_138_0))))) | (i_2_3_86_0 & ((i_2_3_29_0 & ((i_2_3_68_0 & i_2_3_99_0) | (~i_2_3_68_0 & ~i_2_3_99_0 & i_2_3_142_0))) | (i_2_3_68_0 & (~i_2_3_138_0 | (~i_2_3_79_0 & i_2_3_99_0))))))) | (~i_2_3_79_0 & ((~i_2_3_77_0 & ((~i_2_3_43_0 & ~i_2_3_138_0 & (i_2_3_72_0 | i_2_3_99_0)) | (i_2_3_68_0 & ((i_2_3_29_0 & i_2_3_72_0 & i_2_3_99_0) | (~i_2_3_29_0 & ~i_2_3_72_0 & ~i_2_3_86_0 & i_2_3_142_0))) | (i_2_3_29_0 & i_2_3_86_0 & (~i_2_3_72_0 | i_2_3_99_0)))) | (i_2_3_86_0 & ((i_2_3_29_0 & ((i_2_3_68_0 & i_2_3_99_0) | (~i_2_3_43_0 & i_2_3_72_0 & ~i_2_3_99_0))) | (~i_2_3_138_0 & (i_2_3_68_0 | (i_2_3_72_0 & i_2_3_99_0))))) | (i_2_3_43_0 & i_2_3_68_0 & ~i_2_3_138_0))) | (i_2_3_29_0 & ((i_2_3_86_0 & ((i_2_3_99_0 & (~i_2_3_138_0 | (~i_2_3_43_0 & (~i_2_3_77_0 | (i_2_3_68_0 & i_2_3_72_0))))) | (i_2_3_68_0 & ~i_2_3_77_0) | (i_2_3_72_0 & ~i_2_3_138_0))) | (~i_2_3_43_0 & i_2_3_68_0 & ~i_2_3_138_0))) | (~i_2_3_138_0 & ((i_2_3_68_0 & i_2_3_99_0 & (i_2_3_72_0 | ~i_2_3_77_0)) | (~i_2_3_43_0 & ~i_2_3_77_0 & i_2_3_86_0))))) | (i_2_3_68_0 & ((i_2_3_86_0 & ((~i_2_3_77_0 & ((i_2_3_72_0 & ((~i_2_3_79_0 & (~i_2_3_138_0 | (i_2_3_29_0 & (i_2_3_99_0 | ~i_2_3_143_0)))) | (i_2_3_99_0 & ~i_2_3_138_0) | (i_2_3_79_0 & ~i_2_3_143_0 & (i_2_3_99_0 | (~i_2_3_29_0 & ~i_2_3_55_0 & i_2_3_142_0))))) | (~i_2_3_143_0 & ((~i_2_3_79_0 & ~i_2_3_138_0) | (~i_2_3_72_0 & i_2_3_99_0 & (~i_2_3_79_0 | (~i_2_3_29_0 & i_2_3_142_0))))))) | (~i_2_3_43_0 & ~i_2_3_138_0 & ((~i_2_3_79_0 & (i_2_3_99_0 | (i_2_3_72_0 & ~i_2_3_143_0))) | (i_2_3_72_0 & (i_2_3_29_0 | (i_2_3_99_0 & ~i_2_3_143_0))))))) | (~i_2_3_138_0 & ((i_2_3_72_0 & ~i_2_3_77_0 & ((~i_2_3_79_0 & i_2_3_99_0) | (i_2_3_29_0 & ~i_2_3_143_0))) | (i_2_3_29_0 & ((i_2_3_77_0 & (~i_2_3_79_0 | (~i_2_3_72_0 & ~i_2_3_143_0))) | i_2_3_99_0 | (~i_2_3_143_0 & (i_2_3_43_0 | ~i_2_3_79_0)))))))) | (i_2_3_29_0 & ((~i_2_3_138_0 & ((~i_2_3_143_0 & ((~i_2_3_43_0 & i_2_3_99_0 & (i_2_3_72_0 | (i_2_3_77_0 & i_2_3_142_0))) | (~i_2_3_77_0 & i_2_3_86_0) | (~i_2_3_79_0 & (i_2_3_43_0 | i_2_3_77_0)))) | (~i_2_3_77_0 & ((i_2_3_72_0 & ((i_2_3_86_0 & i_2_3_99_0) | (~i_2_3_43_0 & ~i_2_3_79_0))) | (~i_2_3_79_0 & (i_2_3_86_0 | i_2_3_99_0)) | (~i_2_3_72_0 & i_2_3_86_0 & ~i_2_3_99_0))))) | (i_2_3_72_0 & i_2_3_77_0 & ~i_2_3_79_0 & ~i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_143_0))) | (~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_138_0 & ~i_2_3_143_0))) | (i_2_3_29_0 & ((i_2_3_86_0 & ((~i_2_3_43_0 & ((i_2_3_55_0 & i_2_3_68_0 & ~i_2_3_138_0) | (~i_2_3_68_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_143_0))) | (i_2_3_55_0 & ((~i_2_3_77_0 & ((i_2_3_68_0 & (~i_2_3_138_0 | (i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_99_0))) | (~i_2_3_79_0 & (~i_2_3_138_0 | ~i_2_3_143_0)) | (~i_2_3_138_0 & ~i_2_3_143_0) | (i_2_3_99_0 & (~i_2_3_138_0 | (i_2_3_72_0 & ~i_2_3_143_0))))) | (~i_2_3_79_0 & ((i_2_3_99_0 & (~i_2_3_143_0 | (i_2_3_72_0 & ~i_2_3_138_0))) | (i_2_3_68_0 & ~i_2_3_138_0) | (~i_2_3_68_0 & ~i_2_3_143_0))) | (i_2_3_68_0 & ~i_2_3_138_0 & (~i_2_3_72_0 | i_2_3_99_0 | ~i_2_3_143_0)))) | (~i_2_3_138_0 & ((i_2_3_68_0 & ((i_2_3_72_0 & ((~i_2_3_77_0 & (~i_2_3_79_0 | ~i_2_3_143_0)) | (~i_2_3_143_0 & (~i_2_3_79_0 | i_2_3_99_0)))) | (i_2_3_99_0 & (~i_2_3_77_0 | ~i_2_3_79_0)))) | (~i_2_3_77_0 & ~i_2_3_143_0 & (~i_2_3_79_0 | (i_2_3_72_0 & i_2_3_99_0))))))) | (i_2_3_55_0 & ((~i_2_3_77_0 & ((i_2_3_99_0 & ((~i_2_3_43_0 & (~i_2_3_138_0 | (~i_2_3_79_0 & ~i_2_3_143_0))) | (~i_2_3_138_0 & (~i_2_3_79_0 | (i_2_3_68_0 & i_2_3_72_0))))) | (~i_2_3_138_0 & ((i_2_3_68_0 & (~i_2_3_79_0 | (i_2_3_72_0 & ~i_2_3_143_0))) | (i_2_3_72_0 & ~i_2_3_79_0 & ~i_2_3_143_0))))) | (~i_2_3_138_0 & ((i_2_3_68_0 & ~i_2_3_79_0 & i_2_3_99_0) | (~i_2_3_143_0 & ((i_2_3_68_0 & (i_2_3_99_0 | (i_2_3_72_0 & ~i_2_3_79_0))) | (i_2_3_79_0 & i_2_3_99_0 & i_2_3_43_0 & i_2_3_72_0))))))) | (~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_138_0 & ~i_2_3_143_0))) | (i_2_3_55_0 & ((i_2_3_86_0 & ((~i_2_3_138_0 & ((i_2_3_68_0 & (((~i_2_3_77_0 | ~i_2_3_79_0) & (i_2_3_99_0 | (i_2_3_72_0 & ~i_2_3_143_0))) | (~i_2_3_77_0 & ~i_2_3_79_0) | (i_2_3_99_0 & ~i_2_3_143_0))) | (i_2_3_99_0 & ((~i_2_3_72_0 & ~i_2_3_79_0 & (~i_2_3_77_0 | ~i_2_3_143_0)) | (~i_2_3_77_0 & ~i_2_3_143_0))))) | (~i_2_3_43_0 & ~i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & ~i_2_3_143_0))) | (i_2_3_68_0 & ~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_143_0 & ((~i_2_3_77_0 & ~i_2_3_138_0) | (~i_2_3_72_0 & ~i_2_3_86_0 & i_2_3_142_0))))) | (i_2_3_68_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_138_0 & ~i_2_3_143_0))) | (~i_2_3_138_0 & ((i_2_3_29_0 & ((~i_2_3_42_0 & ((i_2_3_86_0 & ((~i_2_3_77_0 & ((~i_2_3_43_0 & ((~i_2_3_79_0 & i_2_3_99_0) | (i_2_3_72_0 & ~i_2_3_99_0 & ~i_2_3_143_0))) | ((~i_2_3_79_0 | i_2_3_99_0) & ((i_2_3_55_0 & i_2_3_72_0) | (i_2_3_68_0 & ~i_2_3_143_0))) | (i_2_3_55_0 & (i_2_3_68_0 | (~i_2_3_79_0 & i_2_3_99_0))) | (i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_79_0))) | (i_2_3_72_0 & ((i_2_3_77_0 & i_2_3_142_0 & ((~i_2_3_79_0 & i_2_3_99_0) | (~i_2_3_68_0 & ~i_2_3_143_0 & (~i_2_3_79_0 | (i_2_3_43_0 & i_2_3_99_0))))) | (i_2_3_55_0 & ((~i_2_3_79_0 & (i_2_3_68_0 | i_2_3_99_0)) | (i_2_3_68_0 & (i_2_3_99_0 | ~i_2_3_143_0)))))) | (i_2_3_55_0 & ~i_2_3_79_0 & ((i_2_3_68_0 & ~i_2_3_143_0) | (i_2_3_43_0 & (i_2_3_68_0 | ~i_2_3_143_0)))))) | (i_2_3_55_0 & ((~i_2_3_77_0 & ((~i_2_3_79_0 & ((~i_2_3_43_0 & ((i_2_3_68_0 & i_2_3_72_0) | (i_2_3_99_0 & ~i_2_3_143_0))) | (i_2_3_68_0 & (i_2_3_99_0 | ~i_2_3_143_0)) | (i_2_3_72_0 & i_2_3_99_0 & ~i_2_3_143_0))) | (i_2_3_68_0 & ((i_2_3_99_0 & ~i_2_3_143_0) | (~i_2_3_43_0 & i_2_3_72_0 & (i_2_3_99_0 | ~i_2_3_143_0)))))) | (~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_143_0 & (i_2_3_68_0 | (i_2_3_43_0 & i_2_3_77_0))))) | (~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_143_0 & i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_77_0))) | (i_2_3_55_0 & ((~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_143_0 & i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_77_0) | (i_2_3_86_0 & ((~i_2_3_143_0 & ((~i_2_3_43_0 & ((i_2_3_68_0 & (~i_2_3_77_0 | (i_2_3_72_0 & ~i_2_3_79_0))) | (i_2_3_72_0 & i_2_3_79_0 & i_2_3_99_0))) | (~i_2_3_79_0 & ((~i_2_3_72_0 & i_2_3_99_0) | (i_2_3_68_0 & (~i_2_3_77_0 | i_2_3_99_0)))))) | (i_2_3_68_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & (~i_2_3_43_0 | i_2_3_99_0)))))) | (i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_143_0))) | (~i_2_3_79_0 & ((i_2_3_86_0 & ((~i_2_3_143_0 & ((~i_2_3_42_0 & ((i_2_3_72_0 & ((i_2_3_43_0 & ((i_2_3_55_0 & ~i_2_3_77_0) | (i_2_3_68_0 & i_2_3_99_0))) | (i_2_3_55_0 & ~i_2_3_77_0 & i_2_3_99_0))) | (i_2_3_55_0 & i_2_3_68_0 & (~i_2_3_77_0 | (~i_2_3_43_0 & i_2_3_99_0))))) | (i_2_3_55_0 & i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_77_0 & i_2_3_99_0))) | (~i_2_3_43_0 & i_2_3_55_0 & i_2_3_68_0 & ~i_2_3_72_0 & ~i_2_3_77_0 & ~i_2_3_99_0))) | (~i_2_3_42_0 & ~i_2_3_43_0 & i_2_3_55_0 & i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_77_0 & i_2_3_99_0 & ~i_2_3_143_0))) | (~i_2_3_42_0 & i_2_3_55_0 & i_2_3_68_0 & ~i_2_3_77_0 & i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_143_0))) | (i_2_3_29_0 & i_2_3_86_0 & ((i_2_3_55_0 & ~i_2_3_77_0 & ((~i_2_3_143_0 & ((i_2_3_72_0 & ((i_2_3_43_0 & i_2_3_79_0 & ((i_2_3_68_0 & i_2_3_99_0) | (~i_2_3_42_0 & ~i_2_3_99_0))) | (~i_2_3_42_0 & ~i_2_3_43_0 & (~i_2_3_79_0 | i_2_3_99_0)))) | (~i_2_3_42_0 & i_2_3_99_0 & ((i_2_3_68_0 & ~i_2_3_79_0) | (~i_2_3_68_0 & i_2_3_79_0 & i_2_3_142_0))))) | (i_2_3_72_0 & ~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_42_0 & ~i_2_3_43_0 & i_2_3_68_0))) | (~i_2_3_42_0 & ~i_2_3_43_0 & i_2_3_72_0 & i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_143_0))))) | (i_2_3_91_0 & ((i_2_3_55_0 & ((i_2_3_86_0 & ((~i_2_3_77_0 & ((~i_2_3_42_0 & ((~i_2_3_43_0 & ((~i_2_3_29_0 & ((i_2_3_72_0 & ~i_2_3_138_0) | (~i_2_3_79_0 & i_2_3_99_0 & i_2_3_142_0 & ~i_2_3_143_0))) | (i_2_3_68_0 & ~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_143_0))) | (i_2_3_142_0 & ((i_2_3_72_0 & ~i_2_3_79_0 & ~i_2_3_138_0) | (i_2_3_29_0 & ~i_2_3_68_0 & ~i_2_3_72_0 & i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_143_0))) | (~i_2_3_79_0 & ((i_2_3_72_0 & ((i_2_3_68_0 & i_2_3_99_0) | (i_2_3_29_0 & ~i_2_3_143_0))) | (i_2_3_68_0 & ~i_2_3_138_0) | (i_2_3_29_0 & ((i_2_3_68_0 & i_2_3_99_0) | (~i_2_3_138_0 & ~i_2_3_143_0))))) | (i_2_3_72_0 & ((i_2_3_68_0 & ~i_2_3_138_0) | (i_2_3_29_0 & i_2_3_43_0 & ~i_2_3_143_0))))) | (~i_2_3_138_0 & ((i_2_3_68_0 & ((i_2_3_72_0 & ((i_2_3_29_0 & (i_2_3_99_0 | ~i_2_3_143_0)) | (~i_2_3_79_0 & (i_2_3_29_0 | (i_2_3_99_0 & ~i_2_3_143_0))))) | (i_2_3_29_0 & ((i_2_3_99_0 & ~i_2_3_143_0) | (~i_2_3_79_0 & (i_2_3_99_0 | ~i_2_3_143_0)))))) | (i_2_3_29_0 & ~i_2_3_79_0 & ~i_2_3_143_0 & (i_2_3_99_0 | (~i_2_3_43_0 & i_2_3_72_0))))))) | (~i_2_3_138_0 & ((~i_2_3_42_0 & ((i_2_3_43_0 & ((i_2_3_68_0 & i_2_3_72_0 & i_2_3_99_0) | (~i_2_3_68_0 & i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_142_0 & ~i_2_3_143_0))) | (i_2_3_68_0 & ((i_2_3_29_0 & (~i_2_3_143_0 | (~i_2_3_43_0 & i_2_3_99_0))) | (i_2_3_99_0 & (~i_2_3_79_0 | (~i_2_3_72_0 & ~i_2_3_143_0))))) | (i_2_3_29_0 & i_2_3_72_0 & ~i_2_3_143_0))) | (i_2_3_29_0 & i_2_3_68_0 & ~i_2_3_143_0 & ((~i_2_3_79_0 & i_2_3_99_0) | (~i_2_3_43_0 & i_2_3_72_0 & (~i_2_3_79_0 | i_2_3_99_0)))))))) | (~i_2_3_138_0 & ((~i_2_3_42_0 & ((~i_2_3_77_0 & ((i_2_3_99_0 & ((i_2_3_68_0 & (i_2_3_29_0 | (i_2_3_72_0 & ~i_2_3_79_0))) | (i_2_3_29_0 & ~i_2_3_79_0 & (~i_2_3_43_0 | i_2_3_143_0)) | (i_2_3_72_0 & i_2_3_79_0 & i_2_3_142_0 & i_2_3_143_0))) | (i_2_3_29_0 & i_2_3_68_0 & (i_2_3_43_0 | (~i_2_3_143_0 & (i_2_3_72_0 | ~i_2_3_79_0)))))) | (~i_2_3_79_0 & i_2_3_143_0 & i_2_3_29_0 & i_2_3_72_0))) | (i_2_3_29_0 & i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_143_0))))) | (~i_2_3_138_0 & ((i_2_3_29_0 & ((i_2_3_68_0 & i_2_3_72_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_143_0) | (~i_2_3_42_0 & ((i_2_3_68_0 & ((i_2_3_72_0 & ((~i_2_3_43_0 & ((i_2_3_77_0 & i_2_3_99_0) | (~i_2_3_77_0 & i_2_3_86_0 & ~i_2_3_143_0))) | (~i_2_3_79_0 & ((~i_2_3_77_0 & i_2_3_143_0) | (i_2_3_77_0 & ~i_2_3_143_0))))) | (~i_2_3_79_0 & i_2_3_99_0) | (~i_2_3_77_0 & i_2_3_86_0 & ~i_2_3_143_0 & (~i_2_3_79_0 | i_2_3_99_0)))) | (~i_2_3_43_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_143_0))))) | (~i_2_3_42_0 & i_2_3_43_0 & i_2_3_68_0 & ~i_2_3_72_0 & ~i_2_3_77_0 & i_2_3_79_0 & ~i_2_3_143_0))))) | (~i_2_3_42_0 & ((i_2_3_86_0 & ((~i_2_3_138_0 & ((~i_2_3_77_0 & ((~i_2_3_79_0 & ((i_2_3_99_0 & ((i_2_3_72_0 & ((i_2_3_29_0 & (~i_2_3_43_0 | (i_2_3_142_0 & ~i_2_3_143_0))) | (i_2_3_68_0 & (i_2_3_55_0 | (~i_2_3_43_0 & i_2_3_142_0))))) | (i_2_3_29_0 & i_2_3_55_0 & i_2_3_68_0))) | (i_2_3_29_0 & ~i_2_3_43_0 & i_2_3_55_0 & i_2_3_68_0 & ~i_2_3_143_0))) | (i_2_3_72_0 & i_2_3_99_0 & ~i_2_3_143_0 & i_2_3_29_0 & i_2_3_68_0))) | (i_2_3_29_0 & i_2_3_55_0 & i_2_3_68_0 & ~i_2_3_72_0 & i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_143_0))) | (i_2_3_29_0 & i_2_3_43_0 & i_2_3_47_0 & i_2_3_55_0 & i_2_3_68_0 & ~i_2_3_79_0 & i_2_3_99_0 & i_2_3_142_0 & ~i_2_3_143_0))) | (i_2_3_55_0 & i_2_3_68_0 & i_2_3_29_0 & ~i_2_3_43_0 & i_2_3_72_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_99_0 & ~i_2_3_138_0))) | (i_2_3_29_0 & ~i_2_3_43_0 & i_2_3_55_0 & i_2_3_72_0 & ~i_2_3_77_0 & ~i_2_3_79_0 & i_2_3_86_0 & i_2_3_99_0 & ~i_2_3_138_0 & ~i_2_3_143_0);
endmodule
