// Benchmark "kernel_2_4" written by ABC on Wed May  4 16:42:57 2022

module kernel_2_4 ( 
    i_2_4_12_0, i_2_4_18_0, i_2_4_22_0, i_2_4_24_0, i_2_4_37_0, i_2_4_42_0,
    i_2_4_57_0, i_2_4_70_0, i_2_4_73_0, i_2_4_94_0, i_2_4_109_0,
    i_2_4_117_0, i_2_4_122_0, i_2_4_123_0, i_2_4_133_0,
    o_2_4_0_0  );
  input  i_2_4_12_0, i_2_4_18_0, i_2_4_22_0, i_2_4_24_0, i_2_4_37_0,
    i_2_4_42_0, i_2_4_57_0, i_2_4_70_0, i_2_4_73_0, i_2_4_94_0,
    i_2_4_109_0, i_2_4_117_0, i_2_4_122_0, i_2_4_123_0, i_2_4_133_0;
  output o_2_4_0_0;
  wire new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_;
  NOT      g000(.a(i_2_4_123_0), .O(new_n17_));
  NOT      g001(.a(i_2_4_133_0), .O(new_n18_));
  NOT      g002(.a(i_2_4_117_0), .O(new_n19_));
  NOT      g003(.a(i_2_4_70_0), .O(new_n20_));
  NOT      g004(.a(i_2_4_42_0), .O(new_n21_));
  OR       g005(.a(i_2_4_122_0), .b(i_2_4_37_0), .O(new_n22_));
  NOT      g006(.a(new_n22_), .O(new_n23_));
  OR       g007(.a(i_2_4_109_0), .b(i_2_4_24_0), .O(new_n24_));
  AND      g008(.a(new_n24_), .b(new_n23_), .O(new_n25_));
  AND      g009(.a(i_2_4_94_0), .b(i_2_4_73_0), .O(new_n26_));
  AND      g010(.a(new_n26_), .b(i_2_4_109_0), .O(new_n27_));
  AND      g011(.a(i_2_4_94_0), .b(i_2_4_24_0), .O(new_n28_));
  OR       g012(.a(new_n28_), .b(new_n27_), .O(new_n29_));
  NOT      g013(.a(i_2_4_37_0), .O(new_n30_));
  AND      g014(.a(i_2_4_73_0), .b(new_n30_), .O(new_n31_));
  NAND     g015(.a(i_2_4_122_0), .b(i_2_4_24_0), .O(new_n32_));
  OR       g016(.a(new_n32_), .b(new_n31_), .O(new_n33_));
  AND      g017(.a(new_n33_), .b(new_n29_), .O(new_n34_));
  OR       g018(.a(new_n34_), .b(new_n25_), .O(new_n35_));
  AND      g019(.a(new_n35_), .b(i_2_4_12_0), .O(new_n36_));
  NOT      g020(.a(i_2_4_122_0), .O(new_n37_));
  AND      g021(.a(new_n37_), .b(i_2_4_73_0), .O(new_n38_));
  AND      g022(.a(new_n37_), .b(i_2_4_24_0), .O(new_n39_));
  OR       g023(.a(new_n39_), .b(i_2_4_18_0), .O(new_n40_));
  AND      g024(.a(new_n40_), .b(i_2_4_109_0), .O(new_n41_));
  OR       g025(.a(new_n41_), .b(new_n38_), .O(new_n42_));
  AND      g026(.a(new_n42_), .b(new_n30_), .O(new_n43_));
  NOT      g027(.a(i_2_4_12_0), .O(new_n44_));
  AND      g028(.a(new_n28_), .b(i_2_4_109_0), .O(new_n45_));
  NOT      g029(.a(new_n24_), .O(new_n46_));
  AND      g030(.a(i_2_4_73_0), .b(i_2_4_18_0), .O(new_n47_));
  AND      g031(.a(new_n47_), .b(new_n46_), .O(new_n48_));
  OR       g032(.a(new_n48_), .b(new_n45_), .O(new_n49_));
  AND      g033(.a(new_n49_), .b(new_n44_), .O(new_n50_));
  OR       g034(.a(new_n50_), .b(new_n43_), .O(new_n51_));
  OR       g035(.a(new_n51_), .b(new_n36_), .O(new_n52_));
  AND      g036(.a(new_n52_), .b(i_2_4_22_0), .O(new_n53_));
  AND      g037(.a(new_n37_), .b(i_2_4_12_0), .O(new_n54_));
  OR       g038(.a(new_n54_), .b(i_2_4_18_0), .O(new_n55_));
  OR       g039(.a(new_n24_), .b(i_2_4_94_0), .O(new_n56_));
  AND      g040(.a(new_n56_), .b(new_n55_), .O(new_n57_));
  AND      g041(.a(i_2_4_109_0), .b(i_2_4_24_0), .O(new_n58_));
  AND      g042(.a(new_n58_), .b(new_n37_), .O(new_n59_));
  OR       g043(.a(new_n59_), .b(new_n57_), .O(new_n60_));
  AND      g044(.a(new_n60_), .b(new_n30_), .O(new_n61_));
  AND      g045(.a(new_n37_), .b(i_2_4_18_0), .O(new_n62_));
  AND      g046(.a(new_n62_), .b(new_n24_), .O(new_n63_));
  OR       g047(.a(new_n63_), .b(new_n61_), .O(new_n64_));
  AND      g048(.a(new_n64_), .b(i_2_4_73_0), .O(new_n65_));
  AND      g049(.a(i_2_4_24_0), .b(i_2_4_12_0), .O(new_n66_));
  AND      g050(.a(new_n66_), .b(i_2_4_109_0), .O(new_n67_));
  OR       g051(.a(new_n67_), .b(new_n30_), .O(new_n68_));
  AND      g052(.a(new_n68_), .b(new_n62_), .O(new_n69_));
  OR       g053(.a(new_n69_), .b(new_n65_), .O(new_n70_));
  OR       g054(.a(new_n70_), .b(new_n53_), .O(new_n71_));
  AND      g055(.a(new_n71_), .b(new_n21_), .O(new_n72_));
  NOT      g056(.a(i_2_4_22_0), .O(new_n73_));
  NOT      g057(.a(i_2_4_94_0), .O(new_n74_));
  NOT      g058(.a(i_2_4_73_0), .O(new_n75_));
  OR       g059(.a(new_n75_), .b(i_2_4_42_0), .O(new_n76_));
  OR       g060(.a(new_n76_), .b(new_n74_), .O(new_n77_));
  NAND     g061(.a(i_2_4_18_0), .b(new_n44_), .O(new_n78_));
  OR       g062(.a(new_n78_), .b(new_n77_), .O(new_n79_));
  AND      g063(.a(new_n30_), .b(i_2_4_24_0), .O(new_n80_));
  AND      g064(.a(new_n75_), .b(i_2_4_42_0), .O(new_n81_));
  AND      g065(.a(new_n81_), .b(new_n54_), .O(new_n82_));
  NAND     g066(.a(new_n82_), .b(new_n80_), .O(new_n83_));
  NAND     g067(.a(new_n83_), .b(new_n79_), .O(new_n84_));
  AND      g068(.a(new_n84_), .b(new_n73_), .O(new_n85_));
  OR       g069(.a(i_2_4_109_0), .b(i_2_4_12_0), .O(new_n86_));
  AND      g070(.a(new_n86_), .b(i_2_4_22_0), .O(new_n87_));
  OR       g071(.a(new_n87_), .b(new_n58_), .O(new_n88_));
  AND      g072(.a(new_n23_), .b(i_2_4_94_0), .O(new_n89_));
  AND      g073(.a(new_n89_), .b(new_n88_), .O(new_n90_));
  OR       g074(.a(new_n90_), .b(new_n85_), .O(new_n91_));
  OR       g075(.a(new_n91_), .b(new_n72_), .O(new_n92_));
  AND      g076(.a(new_n92_), .b(new_n20_), .O(new_n93_));
  OR       g077(.a(i_2_4_94_0), .b(i_2_4_12_0), .O(new_n94_));
  OR       g078(.a(new_n94_), .b(i_2_4_24_0), .O(new_n95_));
  AND      g079(.a(new_n95_), .b(i_2_4_73_0), .O(new_n96_));
  OR       g080(.a(i_2_4_94_0), .b(i_2_4_73_0), .O(new_n97_));
  AND      g081(.a(new_n97_), .b(new_n24_), .O(new_n98_));
  OR       g082(.a(new_n98_), .b(new_n67_), .O(new_n99_));
  OR       g083(.a(new_n99_), .b(new_n96_), .O(new_n100_));
  AND      g084(.a(new_n100_), .b(new_n21_), .O(new_n101_));
  OR       g085(.a(new_n58_), .b(i_2_4_94_0), .O(new_n102_));
  AND      g086(.a(new_n102_), .b(new_n98_), .O(new_n103_));
  AND      g087(.a(new_n103_), .b(i_2_4_12_0), .O(new_n104_));
  OR       g088(.a(new_n104_), .b(new_n45_), .O(new_n105_));
  OR       g089(.a(new_n105_), .b(new_n101_), .O(new_n106_));
  AND      g090(.a(new_n106_), .b(i_2_4_22_0), .O(new_n107_));
  AND      g091(.a(i_2_4_109_0), .b(new_n21_), .O(new_n108_));
  AND      g092(.a(new_n108_), .b(new_n26_), .O(new_n109_));
  AND      g093(.a(i_2_4_109_0), .b(i_2_4_12_0), .O(new_n110_));
  NOT      g094(.a(new_n110_), .O(new_n111_));
  NAND     g095(.a(new_n111_), .b(new_n77_), .O(new_n112_));
  NAND     g096(.a(new_n76_), .b(new_n74_), .O(new_n113_));
  AND      g097(.a(new_n113_), .b(i_2_4_24_0), .O(new_n114_));
  AND      g098(.a(new_n114_), .b(new_n112_), .O(new_n115_));
  OR       g099(.a(new_n115_), .b(new_n109_), .O(new_n116_));
  OR       g100(.a(new_n116_), .b(new_n107_), .O(new_n117_));
  AND      g101(.a(new_n117_), .b(new_n23_), .O(new_n118_));
  AND      g102(.a(new_n21_), .b(i_2_4_22_0), .O(new_n119_));
  AND      g103(.a(new_n119_), .b(i_2_4_24_0), .O(new_n120_));
  AND      g104(.a(i_2_4_94_0), .b(i_2_4_70_0), .O(new_n121_));
  AND      g105(.a(new_n121_), .b(new_n110_), .O(new_n122_));
  AND      g106(.a(new_n122_), .b(new_n120_), .O(new_n123_));
  OR       g107(.a(new_n123_), .b(new_n118_), .O(new_n124_));
  OR       g108(.a(new_n124_), .b(new_n93_), .O(new_n125_));
  AND      g109(.a(new_n125_), .b(new_n19_), .O(new_n126_));
  AND      g110(.a(new_n94_), .b(new_n80_), .O(new_n127_));
  AND      g111(.a(new_n26_), .b(i_2_4_12_0), .O(new_n128_));
  OR       g112(.a(new_n128_), .b(new_n127_), .O(new_n129_));
  AND      g113(.a(new_n129_), .b(i_2_4_109_0), .O(new_n130_));
  OR       g114(.a(new_n110_), .b(i_2_4_22_0), .O(new_n131_));
  OR       g115(.a(new_n131_), .b(i_2_4_73_0), .O(new_n132_));
  NAND     g116(.a(i_2_4_94_0), .b(i_2_4_22_0), .O(new_n133_));
  NAND     g117(.a(new_n133_), .b(i_2_4_37_0), .O(new_n134_));
  AND      g118(.a(new_n134_), .b(new_n132_), .O(new_n135_));
  AND      g119(.a(i_2_4_73_0), .b(i_2_4_12_0), .O(new_n136_));
  AND      g120(.a(new_n136_), .b(new_n24_), .O(new_n137_));
  AND      g121(.a(new_n137_), .b(new_n102_), .O(new_n138_));
  OR       g122(.a(new_n138_), .b(new_n45_), .O(new_n139_));
  OR       g123(.a(new_n139_), .b(i_2_4_22_0), .O(new_n140_));
  AND      g124(.a(new_n140_), .b(i_2_4_24_0), .O(new_n141_));
  OR       g125(.a(new_n141_), .b(new_n135_), .O(new_n142_));
  AND      g126(.a(new_n142_), .b(new_n37_), .O(new_n143_));
  OR       g127(.a(new_n143_), .b(new_n130_), .O(new_n144_));
  AND      g128(.a(new_n144_), .b(new_n20_), .O(new_n145_));
  AND      g129(.a(i_2_4_109_0), .b(i_2_4_73_0), .O(new_n146_));
  OR       g130(.a(new_n146_), .b(new_n80_), .O(new_n147_));
  AND      g131(.a(new_n147_), .b(i_2_4_70_0), .O(new_n148_));
  AND      g132(.a(new_n54_), .b(i_2_4_73_0), .O(new_n149_));
  NAND     g133(.a(i_2_4_122_0), .b(i_2_4_37_0), .O(new_n150_));
  AND      g134(.a(new_n150_), .b(i_2_4_22_0), .O(new_n151_));
  OR       g135(.a(new_n151_), .b(new_n149_), .O(new_n152_));
  OR       g136(.a(new_n152_), .b(new_n148_), .O(new_n153_));
  AND      g137(.a(new_n153_), .b(i_2_4_94_0), .O(new_n154_));
  OR       g138(.a(new_n30_), .b(i_2_4_22_0), .O(new_n155_));
  AND      g139(.a(new_n155_), .b(new_n37_), .O(new_n156_));
  AND      g140(.a(new_n30_), .b(i_2_4_22_0), .O(new_n157_));
  AND      g141(.a(new_n157_), .b(i_2_4_73_0), .O(new_n158_));
  OR       g142(.a(new_n158_), .b(new_n156_), .O(new_n159_));
  AND      g143(.a(new_n159_), .b(i_2_4_109_0), .O(new_n160_));
  OR       g144(.a(i_2_4_24_0), .b(i_2_4_12_0), .O(new_n161_));
  AND      g145(.a(new_n161_), .b(new_n23_), .O(new_n162_));
  OR       g146(.a(new_n162_), .b(new_n160_), .O(new_n163_));
  OR       g147(.a(new_n137_), .b(i_2_4_22_0), .O(new_n164_));
  OR       g148(.a(new_n136_), .b(i_2_4_24_0), .O(new_n165_));
  AND      g149(.a(new_n165_), .b(new_n150_), .O(new_n166_));
  AND      g150(.a(new_n166_), .b(new_n164_), .O(new_n167_));
  NAND     g151(.a(new_n58_), .b(i_2_4_70_0), .O(new_n168_));
  OR       g152(.a(new_n74_), .b(i_2_4_73_0), .O(new_n169_));
  OR       g153(.a(new_n169_), .b(i_2_4_122_0), .O(new_n170_));
  NAND     g154(.a(new_n170_), .b(new_n168_), .O(new_n171_));
  AND      g155(.a(new_n171_), .b(new_n44_), .O(new_n172_));
  OR       g156(.a(new_n172_), .b(new_n167_), .O(new_n173_));
  OR       g157(.a(new_n173_), .b(new_n163_), .O(new_n174_));
  OR       g158(.a(new_n174_), .b(new_n154_), .O(new_n175_));
  AND      g159(.a(new_n175_), .b(new_n21_), .O(new_n176_));
  OR       g160(.a(i_2_4_122_0), .b(i_2_4_24_0), .O(new_n177_));
  AND      g161(.a(new_n177_), .b(i_2_4_12_0), .O(new_n178_));
  OR       g162(.a(new_n178_), .b(new_n156_), .O(new_n179_));
  AND      g163(.a(new_n179_), .b(i_2_4_94_0), .O(new_n180_));
  OR       g164(.a(i_2_4_73_0), .b(i_2_4_24_0), .O(new_n181_));
  AND      g165(.a(new_n181_), .b(new_n23_), .O(new_n182_));
  AND      g166(.a(i_2_4_73_0), .b(i_2_4_24_0), .O(new_n183_));
  AND      g167(.a(i_2_4_42_0), .b(i_2_4_22_0), .O(new_n184_));
  AND      g168(.a(new_n184_), .b(new_n183_), .O(new_n185_));
  OR       g169(.a(new_n185_), .b(new_n182_), .O(new_n186_));
  OR       g170(.a(new_n186_), .b(new_n180_), .O(new_n187_));
  AND      g171(.a(new_n187_), .b(i_2_4_109_0), .O(new_n188_));
  OR       g172(.a(new_n31_), .b(new_n28_), .O(new_n189_));
  AND      g173(.a(new_n189_), .b(i_2_4_22_0), .O(new_n190_));
  AND      g174(.a(new_n95_), .b(new_n31_), .O(new_n191_));
  OR       g175(.a(new_n191_), .b(new_n190_), .O(new_n192_));
  AND      g176(.a(new_n192_), .b(new_n37_), .O(new_n193_));
  OR       g177(.a(new_n193_), .b(new_n188_), .O(new_n194_));
  OR       g178(.a(new_n194_), .b(new_n176_), .O(new_n195_));
  OR       g179(.a(new_n195_), .b(new_n145_), .O(new_n196_));
  AND      g180(.a(new_n196_), .b(new_n19_), .O(new_n197_));
  OR       g181(.a(i_2_4_94_0), .b(new_n20_), .O(new_n198_));
  AND      g182(.a(new_n198_), .b(i_2_4_73_0), .O(new_n199_));
  OR       g183(.a(new_n20_), .b(i_2_4_12_0), .O(new_n200_));
  AND      g184(.a(new_n200_), .b(new_n21_), .O(new_n201_));
  OR       g185(.a(new_n201_), .b(new_n199_), .O(new_n202_));
  AND      g186(.a(new_n202_), .b(new_n30_), .O(new_n203_));
  AND      g187(.a(i_2_4_94_0), .b(new_n21_), .O(new_n204_));
  NAND     g188(.a(i_2_4_73_0), .b(i_2_4_70_0), .O(new_n205_));
  AND      g189(.a(new_n205_), .b(new_n204_), .O(new_n206_));
  OR       g190(.a(new_n206_), .b(new_n203_), .O(new_n207_));
  AND      g191(.a(new_n207_), .b(new_n37_), .O(new_n208_));
  OR       g192(.a(i_2_4_73_0), .b(new_n21_), .O(new_n209_));
  AND      g193(.a(new_n20_), .b(i_2_4_12_0), .O(new_n210_));
  AND      g194(.a(new_n210_), .b(new_n21_), .O(new_n211_));
  OR       g195(.a(new_n211_), .b(new_n37_), .O(new_n212_));
  AND      g196(.a(new_n212_), .b(new_n209_), .O(new_n213_));
  OR       g197(.a(i_2_4_122_0), .b(i_2_4_70_0), .O(new_n214_));
  NAND     g198(.a(new_n214_), .b(new_n76_), .O(new_n215_));
  AND      g199(.a(new_n215_), .b(i_2_4_94_0), .O(new_n216_));
  OR       g200(.a(new_n205_), .b(new_n21_), .O(new_n217_));
  NAND     g201(.a(new_n217_), .b(new_n214_), .O(new_n218_));
  AND      g202(.a(new_n218_), .b(i_2_4_12_0), .O(new_n219_));
  OR       g203(.a(new_n219_), .b(new_n216_), .O(new_n220_));
  OR       g204(.a(new_n220_), .b(new_n213_), .O(new_n221_));
  AND      g205(.a(new_n221_), .b(new_n30_), .O(new_n222_));
  OR       g206(.a(i_2_4_122_0), .b(i_2_4_42_0), .O(new_n223_));
  NOT      g207(.a(new_n223_), .O(new_n224_));
  AND      g208(.a(new_n224_), .b(i_2_4_73_0), .O(new_n225_));
  AND      g209(.a(new_n225_), .b(new_n210_), .O(new_n226_));
  OR       g210(.a(new_n226_), .b(new_n222_), .O(new_n227_));
  AND      g211(.a(new_n227_), .b(i_2_4_109_0), .O(new_n228_));
  OR       g212(.a(new_n228_), .b(new_n208_), .O(new_n229_));
  AND      g213(.a(new_n229_), .b(i_2_4_24_0), .O(new_n230_));
  OR       g214(.a(i_2_4_70_0), .b(i_2_4_12_0), .O(new_n231_));
  OR       g215(.a(new_n231_), .b(new_n74_), .O(new_n232_));
  OR       g216(.a(i_2_4_73_0), .b(new_n20_), .O(new_n233_));
  NAND     g217(.a(new_n233_), .b(new_n54_), .O(new_n234_));
  NAND     g218(.a(new_n234_), .b(new_n232_), .O(new_n235_));
  AND      g219(.a(new_n235_), .b(i_2_4_24_0), .O(new_n236_));
  AND      g220(.a(i_2_4_70_0), .b(new_n30_), .O(new_n237_));
  OR       g221(.a(new_n237_), .b(new_n38_), .O(new_n238_));
  AND      g222(.a(new_n238_), .b(i_2_4_12_0), .O(new_n239_));
  OR       g223(.a(new_n75_), .b(i_2_4_70_0), .O(new_n240_));
  OR       g224(.a(new_n240_), .b(i_2_4_122_0), .O(new_n241_));
  NOT      g225(.a(i_2_4_24_0), .O(new_n242_));
  OR       g226(.a(new_n200_), .b(new_n242_), .O(new_n243_));
  NAND     g227(.a(new_n243_), .b(new_n241_), .O(new_n244_));
  OR       g228(.a(new_n244_), .b(new_n239_), .O(new_n245_));
  AND      g229(.a(new_n245_), .b(new_n21_), .O(new_n246_));
  OR       g230(.a(new_n246_), .b(new_n236_), .O(new_n247_));
  AND      g231(.a(new_n247_), .b(i_2_4_109_0), .O(new_n248_));
  AND      g232(.a(i_2_4_73_0), .b(new_n20_), .O(new_n249_));
  OR       g233(.a(new_n249_), .b(i_2_4_94_0), .O(new_n250_));
  AND      g234(.a(new_n250_), .b(new_n24_), .O(new_n251_));
  AND      g235(.a(i_2_4_94_0), .b(new_n20_), .O(new_n252_));
  OR       g236(.a(new_n252_), .b(new_n37_), .O(new_n253_));
  OR       g237(.a(new_n253_), .b(new_n251_), .O(new_n254_));
  AND      g238(.a(new_n254_), .b(new_n30_), .O(new_n255_));
  OR       g239(.a(new_n250_), .b(new_n183_), .O(new_n256_));
  AND      g240(.a(new_n150_), .b(i_2_4_12_0), .O(new_n257_));
  AND      g241(.a(new_n257_), .b(new_n256_), .O(new_n258_));
  OR       g242(.a(new_n258_), .b(new_n255_), .O(new_n259_));
  AND      g243(.a(new_n259_), .b(new_n21_), .O(new_n260_));
  AND      g244(.a(new_n20_), .b(i_2_4_24_0), .O(new_n261_));
  AND      g245(.a(i_2_4_109_0), .b(new_n44_), .O(new_n262_));
  OR       g246(.a(new_n262_), .b(new_n261_), .O(new_n263_));
  OR       g247(.a(new_n263_), .b(new_n96_), .O(new_n264_));
  AND      g248(.a(new_n264_), .b(new_n23_), .O(new_n265_));
  OR       g249(.a(new_n265_), .b(new_n260_), .O(new_n266_));
  OR       g250(.a(new_n266_), .b(new_n248_), .O(new_n267_));
  AND      g251(.a(new_n267_), .b(i_2_4_22_0), .O(new_n268_));
  OR       g252(.a(new_n268_), .b(new_n230_), .O(new_n269_));
  OR       g253(.a(new_n269_), .b(new_n197_), .O(new_n270_));
  AND      g254(.a(new_n270_), .b(i_2_4_18_0), .O(new_n271_));
  NOT      g255(.a(new_n76_), .O(new_n272_));
  OR       g256(.a(new_n198_), .b(i_2_4_109_0), .O(new_n273_));
  AND      g257(.a(new_n273_), .b(new_n272_), .O(new_n274_));
  AND      g258(.a(new_n200_), .b(i_2_4_94_0), .O(new_n275_));
  OR       g259(.a(new_n275_), .b(new_n211_), .O(new_n276_));
  AND      g260(.a(new_n276_), .b(i_2_4_109_0), .O(new_n277_));
  OR       g261(.a(new_n277_), .b(new_n274_), .O(new_n278_));
  AND      g262(.a(new_n278_), .b(i_2_4_24_0), .O(new_n279_));
  AND      g263(.a(new_n97_), .b(new_n20_), .O(new_n280_));
  AND      g264(.a(new_n280_), .b(new_n112_), .O(new_n281_));
  OR       g265(.a(new_n281_), .b(new_n279_), .O(new_n282_));
  AND      g266(.a(new_n282_), .b(i_2_4_22_0), .O(new_n283_));
  OR       g267(.a(i_2_4_70_0), .b(i_2_4_42_0), .O(new_n284_));
  NOT      g268(.a(new_n284_), .O(new_n285_));
  AND      g269(.a(new_n285_), .b(new_n139_), .O(new_n286_));
  OR       g270(.a(new_n286_), .b(new_n283_), .O(new_n287_));
  AND      g271(.a(new_n287_), .b(new_n30_), .O(new_n288_));
  AND      g272(.a(i_2_4_117_0), .b(i_2_4_70_0), .O(new_n289_));
  AND      g273(.a(new_n289_), .b(new_n27_), .O(new_n290_));
  AND      g274(.a(new_n290_), .b(new_n119_), .O(new_n291_));
  AND      g275(.a(i_2_4_109_0), .b(i_2_4_94_0), .O(new_n292_));
  AND      g276(.a(new_n292_), .b(new_n211_), .O(new_n293_));
  AND      g277(.a(new_n209_), .b(i_2_4_109_0), .O(new_n294_));
  AND      g278(.a(new_n233_), .b(i_2_4_12_0), .O(new_n295_));
  OR       g279(.a(new_n295_), .b(new_n294_), .O(new_n296_));
  AND      g280(.a(new_n296_), .b(i_2_4_94_0), .O(new_n297_));
  OR       g281(.a(i_2_4_109_0), .b(i_2_4_94_0), .O(new_n298_));
  OR       g282(.a(new_n249_), .b(new_n201_), .O(new_n299_));
  AND      g283(.a(new_n299_), .b(new_n298_), .O(new_n300_));
  OR       g284(.a(new_n300_), .b(new_n272_), .O(new_n301_));
  OR       g285(.a(new_n301_), .b(new_n297_), .O(new_n302_));
  AND      g286(.a(new_n302_), .b(new_n30_), .O(new_n303_));
  OR       g287(.a(new_n303_), .b(new_n293_), .O(new_n304_));
  AND      g288(.a(new_n304_), .b(i_2_4_18_0), .O(new_n305_));
  OR       g289(.a(new_n305_), .b(new_n291_), .O(new_n306_));
  OR       g290(.a(new_n306_), .b(new_n288_), .O(new_n307_));
  AND      g291(.a(new_n307_), .b(new_n37_), .O(new_n308_));
  OR       g292(.a(new_n308_), .b(new_n271_), .O(new_n309_));
  OR       g293(.a(new_n309_), .b(new_n126_), .O(new_n310_));
  AND      g294(.a(new_n310_), .b(i_2_4_57_0), .O(new_n311_));
  AND      g295(.a(new_n298_), .b(new_n211_), .O(new_n312_));
  NAND     g296(.a(new_n298_), .b(new_n20_), .O(new_n313_));
  OR       g297(.a(new_n313_), .b(new_n292_), .O(new_n314_));
  NOT      g298(.a(new_n204_), .O(new_n315_));
  NOT      g299(.a(i_2_4_109_0), .O(new_n316_));
  OR       g300(.a(new_n316_), .b(i_2_4_42_0), .O(new_n317_));
  AND      g301(.a(new_n317_), .b(i_2_4_70_0), .O(new_n318_));
  OR       g302(.a(new_n318_), .b(new_n44_), .O(new_n319_));
  AND      g303(.a(new_n319_), .b(new_n315_), .O(new_n320_));
  NAND     g304(.a(new_n320_), .b(new_n314_), .O(new_n321_));
  AND      g305(.a(new_n321_), .b(i_2_4_24_0), .O(new_n322_));
  OR       g306(.a(new_n322_), .b(new_n312_), .O(new_n323_));
  AND      g307(.a(new_n323_), .b(new_n19_), .O(new_n324_));
  AND      g308(.a(new_n24_), .b(new_n20_), .O(new_n325_));
  OR       g309(.a(new_n325_), .b(new_n110_), .O(new_n326_));
  AND      g310(.a(new_n326_), .b(new_n204_), .O(new_n327_));
  OR       g311(.a(new_n327_), .b(new_n324_), .O(new_n328_));
  AND      g312(.a(new_n328_), .b(i_2_4_22_0), .O(new_n329_));
  OR       g313(.a(i_2_4_117_0), .b(i_2_4_70_0), .O(new_n330_));
  NAND     g314(.a(new_n330_), .b(new_n44_), .O(new_n331_));
  AND      g315(.a(new_n204_), .b(new_n58_), .O(new_n332_));
  AND      g316(.a(new_n332_), .b(new_n331_), .O(new_n333_));
  OR       g317(.a(new_n333_), .b(new_n329_), .O(new_n334_));
  AND      g318(.a(new_n334_), .b(i_2_4_73_0), .O(new_n335_));
  AND      g319(.a(new_n66_), .b(i_2_4_22_0), .O(new_n336_));
  AND      g320(.a(new_n252_), .b(new_n19_), .O(new_n337_));
  AND      g321(.a(new_n337_), .b(new_n336_), .O(new_n338_));
  OR       g322(.a(new_n338_), .b(new_n335_), .O(new_n339_));
  AND      g323(.a(new_n339_), .b(new_n23_), .O(new_n340_));
  OR       g324(.a(new_n316_), .b(i_2_4_70_0), .O(new_n341_));
  OR       g325(.a(new_n341_), .b(i_2_4_122_0), .O(new_n342_));
  NAND     g326(.a(new_n237_), .b(new_n316_), .O(new_n343_));
  NAND     g327(.a(new_n343_), .b(new_n342_), .O(new_n344_));
  AND      g328(.a(new_n344_), .b(i_2_4_73_0), .O(new_n345_));
  OR       g329(.a(i_2_4_109_0), .b(new_n20_), .O(new_n346_));
  AND      g330(.a(new_n346_), .b(i_2_4_24_0), .O(new_n347_));
  OR       g331(.a(new_n38_), .b(i_2_4_70_0), .O(new_n348_));
  AND      g332(.a(new_n348_), .b(new_n347_), .O(new_n349_));
  OR       g333(.a(new_n349_), .b(new_n345_), .O(new_n350_));
  AND      g334(.a(new_n350_), .b(i_2_4_94_0), .O(new_n351_));
  AND      g335(.a(i_2_4_109_0), .b(new_n20_), .O(new_n352_));
  OR       g336(.a(new_n352_), .b(i_2_4_73_0), .O(new_n353_));
  AND      g337(.a(new_n353_), .b(new_n30_), .O(new_n354_));
  AND      g338(.a(new_n261_), .b(new_n146_), .O(new_n355_));
  OR       g339(.a(new_n355_), .b(new_n354_), .O(new_n356_));
  AND      g340(.a(new_n356_), .b(new_n37_), .O(new_n357_));
  OR       g341(.a(new_n357_), .b(new_n351_), .O(new_n358_));
  AND      g342(.a(new_n358_), .b(i_2_4_12_0), .O(new_n359_));
  OR       g343(.a(new_n199_), .b(new_n146_), .O(new_n360_));
  OR       g344(.a(i_2_4_94_0), .b(i_2_4_24_0), .O(new_n361_));
  OR       g345(.a(new_n361_), .b(new_n360_), .O(new_n362_));
  OR       g346(.a(new_n346_), .b(i_2_4_73_0), .O(new_n363_));
  AND      g347(.a(new_n363_), .b(new_n37_), .O(new_n364_));
  AND      g348(.a(new_n364_), .b(new_n362_), .O(new_n365_));
  OR       g349(.a(new_n365_), .b(new_n355_), .O(new_n366_));
  AND      g350(.a(new_n366_), .b(new_n30_), .O(new_n367_));
  OR       g351(.a(new_n367_), .b(new_n359_), .O(new_n368_));
  AND      g352(.a(new_n368_), .b(new_n21_), .O(new_n369_));
  NAND     g353(.a(new_n284_), .b(i_2_4_37_0), .O(new_n370_));
  OR       g354(.a(new_n240_), .b(i_2_4_37_0), .O(new_n371_));
  NAND     g355(.a(new_n371_), .b(i_2_4_122_0), .O(new_n372_));
  AND      g356(.a(new_n372_), .b(new_n370_), .O(new_n373_));
  OR       g357(.a(new_n317_), .b(i_2_4_57_0), .O(new_n374_));
  OR       g358(.a(new_n32_), .b(new_n75_), .O(new_n375_));
  NAND     g359(.a(new_n375_), .b(new_n374_), .O(new_n376_));
  AND      g360(.a(new_n376_), .b(new_n44_), .O(new_n377_));
  OR       g361(.a(new_n347_), .b(new_n225_), .O(new_n378_));
  AND      g362(.a(new_n378_), .b(i_2_4_12_0), .O(new_n379_));
  OR       g363(.a(new_n379_), .b(new_n377_), .O(new_n380_));
  OR       g364(.a(new_n380_), .b(new_n373_), .O(new_n381_));
  AND      g365(.a(new_n381_), .b(i_2_4_94_0), .O(new_n382_));
  OR       g366(.a(new_n237_), .b(new_n108_), .O(new_n383_));
  AND      g367(.a(new_n383_), .b(i_2_4_24_0), .O(new_n384_));
  OR       g368(.a(new_n285_), .b(new_n86_), .O(new_n385_));
  AND      g369(.a(new_n385_), .b(new_n30_), .O(new_n386_));
  OR       g370(.a(new_n386_), .b(new_n384_), .O(new_n387_));
  AND      g371(.a(new_n387_), .b(new_n37_), .O(new_n388_));
  OR       g372(.a(i_2_4_70_0), .b(i_2_4_37_0), .O(new_n389_));
  NAND     g373(.a(new_n389_), .b(new_n223_), .O(new_n390_));
  AND      g374(.a(new_n390_), .b(i_2_4_24_0), .O(new_n391_));
  OR       g375(.a(new_n37_), .b(i_2_4_42_0), .O(new_n392_));
  AND      g376(.a(new_n392_), .b(new_n352_), .O(new_n393_));
  OR       g377(.a(new_n393_), .b(new_n391_), .O(new_n394_));
  AND      g378(.a(new_n394_), .b(i_2_4_12_0), .O(new_n395_));
  OR       g379(.a(new_n341_), .b(i_2_4_57_0), .O(new_n396_));
  NAND     g380(.a(new_n396_), .b(new_n223_), .O(new_n397_));
  AND      g381(.a(new_n397_), .b(new_n30_), .O(new_n398_));
  OR       g382(.a(new_n398_), .b(new_n395_), .O(new_n399_));
  AND      g383(.a(new_n399_), .b(i_2_4_73_0), .O(new_n400_));
  OR       g384(.a(new_n400_), .b(new_n388_), .O(new_n401_));
  OR       g385(.a(new_n401_), .b(new_n382_), .O(new_n402_));
  AND      g386(.a(new_n402_), .b(i_2_4_22_0), .O(new_n403_));
  AND      g387(.a(new_n66_), .b(i_2_4_94_0), .O(new_n404_));
  OR       g388(.a(new_n355_), .b(new_n29_), .O(new_n405_));
  AND      g389(.a(new_n405_), .b(new_n37_), .O(new_n406_));
  OR       g390(.a(new_n406_), .b(new_n404_), .O(new_n407_));
  AND      g391(.a(new_n407_), .b(new_n30_), .O(new_n408_));
  OR       g392(.a(new_n408_), .b(new_n403_), .O(new_n409_));
  OR       g393(.a(new_n409_), .b(new_n369_), .O(new_n410_));
  AND      g394(.a(new_n410_), .b(new_n19_), .O(new_n411_));
  AND      g395(.a(new_n298_), .b(new_n200_), .O(new_n412_));
  OR       g396(.a(new_n292_), .b(new_n87_), .O(new_n413_));
  OR       g397(.a(new_n413_), .b(new_n412_), .O(new_n414_));
  AND      g398(.a(new_n414_), .b(i_2_4_73_0), .O(new_n415_));
  OR       g399(.a(new_n110_), .b(i_2_4_94_0), .O(new_n416_));
  NAND     g400(.a(new_n416_), .b(i_2_4_22_0), .O(new_n417_));
  NAND     g401(.a(new_n252_), .b(i_2_4_109_0), .O(new_n418_));
  NAND     g402(.a(new_n418_), .b(new_n417_), .O(new_n419_));
  OR       g403(.a(new_n419_), .b(new_n415_), .O(new_n420_));
  AND      g404(.a(new_n420_), .b(new_n30_), .O(new_n421_));
  AND      g405(.a(new_n313_), .b(new_n44_), .O(new_n422_));
  AND      g406(.a(new_n422_), .b(new_n250_), .O(new_n423_));
  OR       g407(.a(new_n252_), .b(new_n30_), .O(new_n424_));
  AND      g408(.a(new_n424_), .b(i_2_4_12_0), .O(new_n425_));
  OR       g409(.a(new_n425_), .b(new_n31_), .O(new_n426_));
  OR       g410(.a(new_n426_), .b(new_n423_), .O(new_n427_));
  AND      g411(.a(new_n427_), .b(i_2_4_22_0), .O(new_n428_));
  OR       g412(.a(new_n360_), .b(i_2_4_12_0), .O(new_n429_));
  AND      g413(.a(new_n429_), .b(new_n354_), .O(new_n430_));
  OR       g414(.a(new_n430_), .b(new_n290_), .O(new_n431_));
  OR       g415(.a(new_n431_), .b(new_n428_), .O(new_n432_));
  AND      g416(.a(new_n432_), .b(i_2_4_24_0), .O(new_n433_));
  OR       g417(.a(new_n433_), .b(new_n421_), .O(new_n434_));
  AND      g418(.a(new_n434_), .b(new_n21_), .O(new_n435_));
  AND      g419(.a(new_n157_), .b(new_n103_), .O(new_n436_));
  OR       g420(.a(new_n28_), .b(i_2_4_12_0), .O(new_n437_));
  AND      g421(.a(new_n437_), .b(new_n361_), .O(new_n438_));
  OR       g422(.a(new_n438_), .b(new_n131_), .O(new_n439_));
  AND      g423(.a(new_n439_), .b(i_2_4_73_0), .O(new_n440_));
  AND      g424(.a(new_n242_), .b(i_2_4_22_0), .O(new_n441_));
  AND      g425(.a(new_n441_), .b(i_2_4_109_0), .O(new_n442_));
  OR       g426(.a(new_n442_), .b(new_n440_), .O(new_n443_));
  AND      g427(.a(new_n443_), .b(new_n30_), .O(new_n444_));
  AND      g428(.a(new_n146_), .b(new_n74_), .O(new_n445_));
  AND      g429(.a(new_n445_), .b(new_n336_), .O(new_n446_));
  OR       g430(.a(new_n446_), .b(new_n444_), .O(new_n447_));
  AND      g431(.a(new_n447_), .b(new_n20_), .O(new_n448_));
  OR       g432(.a(new_n448_), .b(new_n436_), .O(new_n449_));
  OR       g433(.a(new_n449_), .b(new_n435_), .O(new_n450_));
  AND      g434(.a(new_n450_), .b(new_n37_), .O(new_n451_));
  OR       g435(.a(new_n210_), .b(new_n204_), .O(new_n452_));
  AND      g436(.a(new_n157_), .b(new_n58_), .O(new_n453_));
  AND      g437(.a(new_n453_), .b(new_n452_), .O(new_n454_));
  OR       g438(.a(new_n454_), .b(new_n451_), .O(new_n455_));
  OR       g439(.a(new_n455_), .b(new_n411_), .O(new_n456_));
  AND      g440(.a(new_n456_), .b(i_2_4_18_0), .O(new_n457_));
  OR       g441(.a(new_n457_), .b(new_n340_), .O(new_n458_));
  OR       g442(.a(new_n458_), .b(new_n311_), .O(new_n459_));
  AND      g443(.a(new_n459_), .b(new_n18_), .O(new_n460_));
  AND      g444(.a(new_n20_), .b(i_2_4_57_0), .O(new_n461_));
  NAND     g445(.a(new_n461_), .b(new_n404_), .O(new_n462_));
  OR       g446(.a(new_n19_), .b(i_2_4_57_0), .O(new_n463_));
  NAND     g447(.a(new_n463_), .b(new_n58_), .O(new_n464_));
  NAND     g448(.a(i_2_4_109_0), .b(i_2_4_57_0), .O(new_n465_));
  AND      g449(.a(new_n465_), .b(new_n330_), .O(new_n466_));
  NOT      g450(.a(new_n466_), .O(new_n467_));
  OR       g451(.a(new_n467_), .b(new_n464_), .O(new_n468_));
  OR       g452(.a(new_n468_), .b(new_n319_), .O(new_n469_));
  NAND     g453(.a(new_n469_), .b(new_n462_), .O(new_n470_));
  AND      g454(.a(new_n470_), .b(i_2_4_22_0), .O(new_n471_));
  AND      g455(.a(new_n438_), .b(new_n346_), .O(new_n472_));
  AND      g456(.a(new_n352_), .b(new_n95_), .O(new_n473_));
  OR       g457(.a(new_n473_), .b(new_n472_), .O(new_n474_));
  AND      g458(.a(new_n474_), .b(new_n19_), .O(new_n475_));
  AND      g459(.a(new_n292_), .b(new_n261_), .O(new_n476_));
  OR       g460(.a(new_n476_), .b(new_n475_), .O(new_n477_));
  AND      g461(.a(new_n477_), .b(new_n21_), .O(new_n478_));
  AND      g462(.a(new_n45_), .b(i_2_4_12_0), .O(new_n479_));
  OR       g463(.a(new_n479_), .b(new_n478_), .O(new_n480_));
  AND      g464(.a(new_n480_), .b(i_2_4_73_0), .O(new_n481_));
  AND      g465(.a(new_n337_), .b(new_n67_), .O(new_n482_));
  OR       g466(.a(new_n482_), .b(new_n481_), .O(new_n483_));
  AND      g467(.a(new_n483_), .b(i_2_4_57_0), .O(new_n484_));
  NAND     g468(.a(new_n26_), .b(i_2_4_109_0), .O(new_n485_));
  NAND     g469(.a(new_n330_), .b(new_n485_), .O(new_n486_));
  NAND     g470(.a(i_2_4_73_0), .b(i_2_4_57_0), .O(new_n487_));
  NAND     g471(.a(new_n487_), .b(new_n465_), .O(new_n488_));
  AND      g472(.a(new_n488_), .b(new_n486_), .O(new_n489_));
  AND      g473(.a(new_n19_), .b(i_2_4_57_0), .O(new_n490_));
  OR       g474(.a(new_n490_), .b(new_n121_), .O(new_n491_));
  AND      g475(.a(new_n491_), .b(i_2_4_24_0), .O(new_n492_));
  OR       g476(.a(new_n492_), .b(new_n337_), .O(new_n493_));
  OR       g477(.a(new_n493_), .b(new_n489_), .O(new_n494_));
  AND      g478(.a(new_n494_), .b(i_2_4_12_0), .O(new_n495_));
  NAND     g479(.a(new_n490_), .b(i_2_4_73_0), .O(new_n496_));
  NAND     g480(.a(new_n496_), .b(new_n232_), .O(new_n497_));
  AND      g481(.a(new_n497_), .b(new_n24_), .O(new_n498_));
  OR       g482(.a(new_n487_), .b(new_n289_), .O(new_n499_));
  NAND     g483(.a(new_n499_), .b(new_n464_), .O(new_n500_));
  AND      g484(.a(new_n500_), .b(i_2_4_94_0), .O(new_n501_));
  OR       g485(.a(new_n501_), .b(new_n498_), .O(new_n502_));
  OR       g486(.a(new_n502_), .b(new_n495_), .O(new_n503_));
  AND      g487(.a(new_n503_), .b(new_n21_), .O(new_n504_));
  OR       g488(.a(new_n466_), .b(new_n44_), .O(new_n505_));
  OR       g489(.a(new_n341_), .b(new_n94_), .O(new_n506_));
  NAND     g490(.a(new_n506_), .b(new_n505_), .O(new_n507_));
  AND      g491(.a(new_n507_), .b(i_2_4_73_0), .O(new_n508_));
  AND      g492(.a(new_n19_), .b(i_2_4_109_0), .O(new_n509_));
  AND      g493(.a(new_n509_), .b(new_n198_), .O(new_n510_));
  OR       g494(.a(new_n510_), .b(new_n252_), .O(new_n511_));
  AND      g495(.a(new_n511_), .b(i_2_4_57_0), .O(new_n512_));
  OR       g496(.a(new_n512_), .b(new_n508_), .O(new_n513_));
  AND      g497(.a(new_n513_), .b(i_2_4_24_0), .O(new_n514_));
  AND      g498(.a(new_n19_), .b(i_2_4_94_0), .O(new_n515_));
  NOT      g499(.a(new_n515_), .O(new_n516_));
  OR       g500(.a(new_n499_), .b(new_n19_), .O(new_n517_));
  NAND     g501(.a(new_n517_), .b(new_n516_), .O(new_n518_));
  AND      g502(.a(new_n518_), .b(i_2_4_12_0), .O(new_n519_));
  AND      g503(.a(new_n337_), .b(i_2_4_57_0), .O(new_n520_));
  OR       g504(.a(new_n520_), .b(new_n519_), .O(new_n521_));
  AND      g505(.a(new_n521_), .b(i_2_4_109_0), .O(new_n522_));
  OR       g506(.a(new_n522_), .b(new_n514_), .O(new_n523_));
  OR       g507(.a(new_n523_), .b(new_n504_), .O(new_n524_));
  AND      g508(.a(new_n524_), .b(i_2_4_22_0), .O(new_n525_));
  AND      g509(.a(new_n515_), .b(i_2_4_73_0), .O(new_n526_));
  AND      g510(.a(new_n526_), .b(new_n67_), .O(new_n527_));
  OR       g511(.a(new_n527_), .b(new_n525_), .O(new_n528_));
  OR       g512(.a(new_n528_), .b(new_n484_), .O(new_n529_));
  AND      g513(.a(new_n529_), .b(new_n37_), .O(new_n530_));
  OR       g514(.a(new_n530_), .b(new_n471_), .O(new_n531_));
  AND      g515(.a(new_n531_), .b(new_n30_), .O(new_n532_));
  AND      g516(.a(new_n292_), .b(new_n19_), .O(new_n533_));
  AND      g517(.a(new_n533_), .b(new_n461_), .O(new_n534_));
  AND      g518(.a(new_n534_), .b(new_n120_), .O(new_n535_));
  OR       g519(.a(new_n535_), .b(new_n532_), .O(new_n536_));
  AND      g520(.a(new_n536_), .b(i_2_4_18_0), .O(new_n537_));
  AND      g521(.a(new_n204_), .b(new_n31_), .O(new_n538_));
  AND      g522(.a(new_n538_), .b(new_n490_), .O(new_n539_));
  NOT      g523(.a(new_n342_), .O(new_n540_));
  AND      g524(.a(new_n540_), .b(new_n336_), .O(new_n541_));
  AND      g525(.a(new_n541_), .b(new_n539_), .O(new_n542_));
  OR       g526(.a(new_n542_), .b(new_n537_), .O(new_n543_));
  OR       g527(.a(new_n543_), .b(new_n460_), .O(new_n544_));
  AND      g528(.a(new_n544_), .b(new_n17_), .O(new_n545_));
  AND      g529(.a(new_n18_), .b(i_2_4_73_0), .O(new_n546_));
  NAND     g530(.a(new_n546_), .b(new_n108_), .O(new_n547_));
  OR       g531(.a(new_n18_), .b(i_2_4_22_0), .O(new_n548_));
  OR       g532(.a(new_n548_), .b(new_n343_), .O(new_n549_));
  NAND     g533(.a(new_n549_), .b(new_n547_), .O(new_n550_));
  AND      g534(.a(new_n550_), .b(new_n515_), .O(new_n551_));
  AND      g535(.a(new_n252_), .b(i_2_4_117_0), .O(new_n552_));
  OR       g536(.a(new_n31_), .b(i_2_4_94_0), .O(new_n553_));
  OR       g537(.a(new_n26_), .b(new_n19_), .O(new_n554_));
  AND      g538(.a(new_n554_), .b(new_n18_), .O(new_n555_));
  AND      g539(.a(new_n555_), .b(new_n553_), .O(new_n556_));
  OR       g540(.a(new_n556_), .b(new_n316_), .O(new_n557_));
  NAND     g541(.a(new_n371_), .b(new_n316_), .O(new_n558_));
  AND      g542(.a(new_n558_), .b(new_n21_), .O(new_n559_));
  AND      g543(.a(new_n559_), .b(new_n557_), .O(new_n560_));
  OR       g544(.a(new_n560_), .b(new_n552_), .O(new_n561_));
  AND      g545(.a(new_n561_), .b(i_2_4_22_0), .O(new_n562_));
  OR       g546(.a(new_n562_), .b(new_n551_), .O(new_n563_));
  AND      g547(.a(new_n563_), .b(i_2_4_57_0), .O(new_n564_));
  NOT      g548(.a(new_n418_), .O(new_n565_));
  AND      g549(.a(new_n565_), .b(new_n158_), .O(new_n566_));
  OR       g550(.a(new_n566_), .b(new_n564_), .O(new_n567_));
  AND      g551(.a(new_n567_), .b(i_2_4_12_0), .O(new_n568_));
  AND      g552(.a(new_n113_), .b(new_n44_), .O(new_n569_));
  OR       g553(.a(new_n569_), .b(i_2_4_117_0), .O(new_n570_));
  OR       g554(.a(new_n204_), .b(new_n19_), .O(new_n571_));
  AND      g555(.a(new_n571_), .b(new_n352_), .O(new_n572_));
  AND      g556(.a(new_n572_), .b(new_n570_), .O(new_n573_));
  OR       g557(.a(new_n573_), .b(new_n539_), .O(new_n574_));
  AND      g558(.a(new_n574_), .b(i_2_4_22_0), .O(new_n575_));
  NOT      g559(.a(new_n231_), .O(new_n576_));
  AND      g560(.a(new_n576_), .b(new_n272_), .O(new_n577_));
  AND      g561(.a(new_n577_), .b(new_n533_), .O(new_n578_));
  OR       g562(.a(new_n578_), .b(new_n575_), .O(new_n579_));
  AND      g563(.a(new_n579_), .b(new_n18_), .O(new_n580_));
  OR       g564(.a(new_n580_), .b(new_n568_), .O(new_n581_));
  AND      g565(.a(new_n581_), .b(i_2_4_24_0), .O(new_n582_));
  AND      g566(.a(new_n552_), .b(i_2_4_109_0), .O(new_n583_));
  AND      g567(.a(new_n424_), .b(new_n19_), .O(new_n584_));
  AND      g568(.a(new_n584_), .b(new_n512_), .O(new_n585_));
  OR       g569(.a(new_n585_), .b(new_n583_), .O(new_n586_));
  AND      g570(.a(new_n586_), .b(i_2_4_12_0), .O(new_n587_));
  OR       g571(.a(new_n587_), .b(new_n534_), .O(new_n588_));
  AND      g572(.a(new_n546_), .b(new_n119_), .O(new_n589_));
  AND      g573(.a(new_n589_), .b(new_n588_), .O(new_n590_));
  OR       g574(.a(new_n590_), .b(new_n582_), .O(new_n591_));
  AND      g575(.a(new_n591_), .b(new_n62_), .O(new_n592_));
  OR       g576(.a(new_n592_), .b(new_n545_), .O(o_2_4_0_0));
endmodule


