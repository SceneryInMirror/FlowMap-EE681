module kernel_2_1 ( 
    i_2_1_13_0, i_2_1_32_0, i_2_1_34_0, i_2_1_38_0, i_2_1_41_0, i_2_1_46_0,
    i_2_1_47_0, i_2_1_49_0, i_2_1_51_0, i_2_1_54_0, i_2_1_57_0, i_2_1_68_0,
    i_2_1_70_0, i_2_1_135_0, i_2_1_136_0,
    o_2_1_0_0  );
  input  i_2_1_13_0, i_2_1_32_0, i_2_1_34_0, i_2_1_38_0, i_2_1_41_0,
    i_2_1_46_0, i_2_1_47_0, i_2_1_49_0, i_2_1_51_0, i_2_1_54_0, i_2_1_57_0,
    i_2_1_68_0, i_2_1_70_0, i_2_1_135_0, i_2_1_136_0;
  output o_2_1_0_0;
  assign o_2_1_0_0 = (~i_2_1_47_0 & ((~i_2_1_51_0 & ((~i_2_1_13_0 & ((i_2_1_38_0 & i_2_1_41_0 & ~i_2_1_54_0 & i_2_1_68_0) | (i_2_1_32_0 & i_2_1_34_0 & ~i_2_1_49_0 & ~i_2_1_57_0 & ~i_2_1_135_0 & ~i_2_1_136_0))) | (((i_2_1_38_0 & ~i_2_1_46_0 & i_2_1_135_0) | (i_2_1_70_0 & i_2_1_136_0)) & ((i_2_1_32_0 & i_2_1_34_0 & ~i_2_1_54_0) | (i_2_1_13_0 & ~i_2_1_32_0 & ~i_2_1_57_0))) | (i_2_1_32_0 & ((~i_2_1_46_0 & ((i_2_1_41_0 & ((i_2_1_13_0 & (~i_2_1_57_0 | (i_2_1_68_0 & i_2_1_136_0))) | (~i_2_1_54_0 & ((i_2_1_34_0 & i_2_1_70_0) | (~i_2_1_49_0 & ~i_2_1_70_0))) | (i_2_1_34_0 & ((~i_2_1_49_0 & i_2_1_70_0) | (~i_2_1_70_0 & i_2_1_135_0 & ~i_2_1_136_0))) | (~i_2_1_49_0 & ((~i_2_1_57_0 & (i_2_1_68_0 | (~i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_68_0 & (i_2_1_70_0 | (i_2_1_135_0 & i_2_1_136_0))))) | (i_2_1_135_0 & ((~i_2_1_57_0 & i_2_1_136_0 & (i_2_1_68_0 | i_2_1_70_0)) | (i_2_1_70_0 & (i_2_1_38_0 | i_2_1_68_0)))) | (i_2_1_68_0 & i_2_1_70_0 & i_2_1_136_0))) | (i_2_1_13_0 & ((i_2_1_34_0 & (~i_2_1_54_0 | i_2_1_68_0)) | (i_2_1_38_0 & (~i_2_1_49_0 | (i_2_1_68_0 & i_2_1_135_0))) | (i_2_1_68_0 & (((~i_2_1_49_0 | i_2_1_135_0) & (~i_2_1_57_0 | i_2_1_70_0)) | (i_2_1_135_0 & (~i_2_1_49_0 | i_2_1_136_0)) | ~i_2_1_54_0 | (~i_2_1_57_0 & i_2_1_136_0))))) | (~i_2_1_49_0 & (((~i_2_1_54_0 | i_2_1_68_0) & ((i_2_1_38_0 & i_2_1_70_0) | (i_2_1_34_0 & i_2_1_135_0))) | ((i_2_1_38_0 | i_2_1_70_0) & ((i_2_1_34_0 & ~i_2_1_54_0) | (i_2_1_68_0 & (~i_2_1_57_0 | i_2_1_135_0 | i_2_1_136_0)))) | (~i_2_1_57_0 & (~i_2_1_54_0 | (i_2_1_68_0 & i_2_1_135_0 & i_2_1_136_0))) | (~i_2_1_54_0 & i_2_1_68_0 & (i_2_1_70_0 | i_2_1_135_0)) | (i_2_1_38_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_34_0 & ((~i_2_1_57_0 & (i_2_1_136_0 | (~i_2_1_54_0 & i_2_1_135_0))) | (i_2_1_70_0 & (i_2_1_68_0 | (~i_2_1_54_0 & i_2_1_135_0))) | (i_2_1_68_0 & i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_54_0 & (i_2_1_68_0 | (i_2_1_135_0 & i_2_1_136_0))))) | (i_2_1_68_0 & ((~i_2_1_54_0 & (~i_2_1_57_0 | (i_2_1_135_0 & i_2_1_136_0))) | (~i_2_1_57_0 & i_2_1_70_0 & (i_2_1_135_0 | i_2_1_136_0)))) | (i_2_1_38_0 & ~i_2_1_57_0 & i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_41_0 & ((i_2_1_49_0 & ((i_2_1_57_0 & ((~i_2_1_54_0 & ~i_2_1_135_0 & i_2_1_136_0) | (i_2_1_135_0 & ~i_2_1_136_0 & i_2_1_13_0 & i_2_1_68_0))) | (~i_2_1_57_0 & i_2_1_68_0 & i_2_1_70_0))) | (i_2_1_135_0 & ((~i_2_1_57_0 & ((i_2_1_13_0 & ((i_2_1_68_0 & i_2_1_136_0) | (~i_2_1_49_0 & ~i_2_1_136_0))) | (i_2_1_38_0 & (~i_2_1_54_0 | (~i_2_1_34_0 & i_2_1_46_0 & ~i_2_1_136_0))) | (~i_2_1_54_0 & (i_2_1_34_0 | i_2_1_68_0)) | (i_2_1_68_0 & (i_2_1_70_0 | (~i_2_1_49_0 & i_2_1_136_0))))) | (i_2_1_136_0 & ((i_2_1_34_0 & i_2_1_70_0) | (~i_2_1_49_0 & ((i_2_1_34_0 & (~i_2_1_54_0 | i_2_1_68_0)) | (i_2_1_68_0 & (i_2_1_13_0 | i_2_1_38_0 | ~i_2_1_54_0 | i_2_1_70_0)))))))) | (i_2_1_13_0 & ((i_2_1_38_0 & (~i_2_1_49_0 | ~i_2_1_57_0)) | (~i_2_1_49_0 & ((i_2_1_68_0 & i_2_1_70_0) | (~i_2_1_57_0 & ~i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_68_0 & (i_2_1_34_0 | ~i_2_1_54_0)))) | (i_2_1_38_0 & ((i_2_1_34_0 & ~i_2_1_49_0) | (~i_2_1_57_0 & i_2_1_68_0 & i_2_1_136_0))) | (i_2_1_70_0 & ((i_2_1_34_0 & ~i_2_1_49_0 & (~i_2_1_54_0 | i_2_1_68_0)) | (~i_2_1_57_0 & i_2_1_68_0 & i_2_1_136_0) | (~i_2_1_54_0 & (i_2_1_68_0 | i_2_1_136_0)))) | (~i_2_1_54_0 & ((i_2_1_34_0 & ((~i_2_1_49_0 & i_2_1_68_0) | (~i_2_1_57_0 & ~i_2_1_136_0))) | (~i_2_1_49_0 & ~i_2_1_57_0 & i_2_1_68_0))))) | (~i_2_1_57_0 & ((i_2_1_49_0 & ((i_2_1_38_0 & ~i_2_1_54_0 & i_2_1_70_0) | (i_2_1_34_0 & i_2_1_68_0 & i_2_1_136_0))) | (i_2_1_38_0 & ((~i_2_1_54_0 & ((~i_2_1_49_0 & i_2_1_68_0) | (i_2_1_34_0 & i_2_1_136_0))) | (i_2_1_34_0 & (i_2_1_70_0 | (~i_2_1_41_0 & i_2_1_135_0))) | (~i_2_1_49_0 & (i_2_1_13_0 | (i_2_1_68_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_13_0 & ((i_2_1_68_0 & i_2_1_135_0) | (~i_2_1_68_0 & ~i_2_1_135_0))) | (i_2_1_68_0 & i_2_1_70_0 & ~i_2_1_135_0))) | (~i_2_1_54_0 & ((i_2_1_34_0 & (i_2_1_68_0 | i_2_1_70_0)) | (~i_2_1_49_0 & (i_2_1_13_0 | (~i_2_1_41_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_13_0 & (i_2_1_70_0 | (i_2_1_68_0 & i_2_1_136_0))))) | (i_2_1_13_0 & ((i_2_1_68_0 & i_2_1_70_0) | (i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_41_0 & ~i_2_1_49_0))) | (~i_2_1_49_0 & ((i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_41_0 & i_2_1_70_0) | (~i_2_1_135_0 & ~i_2_1_136_0 & i_2_1_34_0 & i_2_1_68_0))))) | (i_2_1_68_0 & ((i_2_1_136_0 & ((~i_2_1_54_0 & ((i_2_1_34_0 & i_2_1_135_0) | (~i_2_1_41_0 & ~i_2_1_49_0 & i_2_1_57_0 & ~i_2_1_135_0))) | (i_2_1_13_0 & i_2_1_70_0 & ~i_2_1_135_0))) | (~i_2_1_54_0 & (((i_2_1_13_0 | i_2_1_38_0) & (i_2_1_34_0 | i_2_1_70_0)) | (i_2_1_135_0 & (i_2_1_38_0 | i_2_1_70_0 | (i_2_1_34_0 & ~i_2_1_49_0))))) | (i_2_1_38_0 & ~i_2_1_49_0 & i_2_1_135_0 & (i_2_1_13_0 | i_2_1_34_0)))) | (i_2_1_13_0 & (((~i_2_1_49_0 | i_2_1_70_0) & ((i_2_1_34_0 & i_2_1_135_0) | (i_2_1_38_0 & i_2_1_136_0))) | (~i_2_1_49_0 & ((~i_2_1_54_0 & i_2_1_135_0) | (i_2_1_38_0 & (~i_2_1_54_0 | i_2_1_70_0)))))) | (i_2_1_70_0 & i_2_1_136_0 & ((i_2_1_34_0 & (i_2_1_38_0 | (~i_2_1_49_0 & i_2_1_135_0))) | (~i_2_1_49_0 & ~i_2_1_54_0 & i_2_1_135_0))))) | (i_2_1_68_0 & ((i_2_1_34_0 & ((~i_2_1_41_0 & ((i_2_1_13_0 & i_2_1_136_0) | (~i_2_1_57_0 & ~i_2_1_135_0 & ~i_2_1_136_0 & i_2_1_49_0 & ~i_2_1_54_0))) | ((i_2_1_13_0 | ~i_2_1_54_0) & ((~i_2_1_46_0 & ~i_2_1_49_0) | (i_2_1_38_0 & ~i_2_1_57_0) | (i_2_1_49_0 & i_2_1_70_0))) | (~i_2_1_46_0 & ((i_2_1_13_0 & (~i_2_1_54_0 | ~i_2_1_57_0)) | ((~i_2_1_54_0 | i_2_1_135_0) & (i_2_1_38_0 | i_2_1_41_0)) | ((i_2_1_135_0 | i_2_1_136_0) & (~i_2_1_54_0 | (~i_2_1_49_0 & i_2_1_70_0))) | (i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_49_0 & ((i_2_1_135_0 & i_2_1_136_0) | (i_2_1_41_0 & i_2_1_70_0))))) | (i_2_1_13_0 & ((i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_49_0 & ~i_2_1_54_0))) | (~i_2_1_57_0 & ((i_2_1_41_0 & ~i_2_1_49_0) | (~i_2_1_54_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_41_0 & ((~i_2_1_49_0 & i_2_1_136_0 & (~i_2_1_54_0 | i_2_1_70_0)) | (~i_2_1_54_0 & (i_2_1_70_0 | i_2_1_135_0)) | (i_2_1_70_0 & i_2_1_135_0 & ~i_2_1_136_0))) | (~i_2_1_54_0 & i_2_1_135_0 & (i_2_1_70_0 | (~i_2_1_49_0 & i_2_1_136_0))) | (i_2_1_38_0 & i_2_1_49_0 & i_2_1_136_0))) | (~i_2_1_54_0 & ((i_2_1_38_0 & ((~i_2_1_57_0 & i_2_1_136_0) | (i_2_1_13_0 & ~i_2_1_46_0))) | ((~i_2_1_57_0 | i_2_1_70_0) & ((~i_2_1_46_0 & (i_2_1_13_0 | (i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_135_0 & i_2_1_136_0 & i_2_1_41_0 & ~i_2_1_49_0))) | ((i_2_1_70_0 | i_2_1_135_0) & ((~i_2_1_46_0 & ~i_2_1_49_0 & (~i_2_1_57_0 | i_2_1_136_0)) | (i_2_1_13_0 & i_2_1_41_0))) | (i_2_1_135_0 & ((~i_2_1_46_0 & ((i_2_1_13_0 & (~i_2_1_49_0 | i_2_1_136_0)) | (i_2_1_41_0 & (i_2_1_70_0 | i_2_1_136_0)))) | (i_2_1_13_0 & ~i_2_1_49_0 & i_2_1_136_0))))) | (i_2_1_13_0 & ((i_2_1_41_0 & ((i_2_1_38_0 & (~i_2_1_57_0 | (~i_2_1_49_0 & i_2_1_136_0))) | (~i_2_1_46_0 & (((~i_2_1_49_0 | i_2_1_136_0) & (i_2_1_70_0 | i_2_1_135_0)) | (i_2_1_70_0 & i_2_1_135_0))) | (~i_2_1_49_0 & i_2_1_135_0 & i_2_1_136_0 & (~i_2_1_57_0 | i_2_1_70_0)))) | (~i_2_1_46_0 & ((i_2_1_38_0 & (i_2_1_70_0 | (i_2_1_135_0 & i_2_1_136_0))) | ((~i_2_1_57_0 | i_2_1_70_0) & ((i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_49_0 & (i_2_1_135_0 | i_2_1_136_0)))) | (~i_2_1_49_0 & ~i_2_1_57_0 & i_2_1_70_0))) | (i_2_1_38_0 & i_2_1_135_0 & (i_2_1_70_0 | (~i_2_1_49_0 & ~i_2_1_57_0))))) | (i_2_1_38_0 & ((~i_2_1_46_0 & ((i_2_1_41_0 & ((~i_2_1_49_0 & i_2_1_136_0) | (i_2_1_49_0 & i_2_1_135_0 & ~i_2_1_136_0))) | (i_2_1_70_0 & ((~i_2_1_49_0 & (~i_2_1_57_0 | i_2_1_135_0)) | (~i_2_1_57_0 & i_2_1_135_0))))) | (i_2_1_136_0 & ((~i_2_1_49_0 & (i_2_1_70_0 | (i_2_1_41_0 & ~i_2_1_57_0 & i_2_1_135_0))) | (i_2_1_70_0 & (i_2_1_46_0 | i_2_1_135_0)))))) | (~i_2_1_49_0 & ((i_2_1_41_0 & ((~i_2_1_46_0 & ((i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_57_0 & (i_2_1_70_0 | (i_2_1_135_0 & i_2_1_136_0))))) | (i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_57_0 & i_2_1_70_0))) | (i_2_1_70_0 & i_2_1_136_0 & ~i_2_1_46_0 & ~i_2_1_57_0))))) | (i_2_1_38_0 & ((i_2_1_46_0 & ((i_2_1_13_0 & i_2_1_34_0 & i_2_1_49_0 & i_2_1_54_0) | (~i_2_1_54_0 & i_2_1_70_0 & i_2_1_135_0))) | (~i_2_1_49_0 & ((i_2_1_13_0 & ((i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_54_0 & ~i_2_1_57_0))) | (i_2_1_34_0 & ((~i_2_1_54_0 & i_2_1_135_0) | (~i_2_1_46_0 & i_2_1_70_0))) | (i_2_1_54_0 & ((~i_2_1_46_0 & ~i_2_1_57_0 & i_2_1_136_0) | (i_2_1_41_0 & i_2_1_57_0 & i_2_1_70_0 & ~i_2_1_136_0))) | (~i_2_1_54_0 & ((i_2_1_70_0 & i_2_1_135_0) | (~i_2_1_57_0 & ((~i_2_1_46_0 & i_2_1_70_0) | (i_2_1_41_0 & i_2_1_136_0))))) | (i_2_1_41_0 & ~i_2_1_46_0 & (i_2_1_70_0 | ~i_2_1_135_0)))) | (~i_2_1_46_0 & ((i_2_1_13_0 & ((i_2_1_34_0 & ~i_2_1_54_0) | (i_2_1_41_0 & i_2_1_70_0 & i_2_1_136_0))) | (i_2_1_34_0 & (i_2_1_41_0 | (~i_2_1_54_0 & i_2_1_70_0))) | (~i_2_1_57_0 & ((~i_2_1_54_0 & i_2_1_135_0) | (i_2_1_41_0 & i_2_1_136_0))) | (~i_2_1_54_0 & i_2_1_136_0 & (i_2_1_49_0 | i_2_1_70_0)))) | (i_2_1_34_0 & ((i_2_1_13_0 & (i_2_1_41_0 | i_2_1_135_0)) | (i_2_1_41_0 & i_2_1_70_0) | (~i_2_1_57_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_13_0 & ((~i_2_1_57_0 & ~i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_54_0 & (i_2_1_136_0 | (i_2_1_70_0 & i_2_1_135_0))))))) | (~i_2_1_57_0 & ((~i_2_1_135_0 & ((i_2_1_13_0 & i_2_1_41_0 & ~i_2_1_54_0) | (i_2_1_34_0 & i_2_1_70_0 & i_2_1_136_0))) | (~i_2_1_54_0 & ((i_2_1_13_0 & ((~i_2_1_49_0 & i_2_1_135_0) | (i_2_1_41_0 & i_2_1_136_0))) | (i_2_1_41_0 & (~i_2_1_46_0 | i_2_1_70_0)) | (i_2_1_70_0 & ((~i_2_1_49_0 & i_2_1_136_0) | (i_2_1_34_0 & ~i_2_1_46_0 & i_2_1_135_0))) | (~i_2_1_49_0 & ((i_2_1_34_0 & (~i_2_1_46_0 | i_2_1_135_0)) | (~i_2_1_38_0 & ~i_2_1_46_0 & i_2_1_136_0))))) | (i_2_1_13_0 & ((i_2_1_34_0 & i_2_1_135_0) | (i_2_1_70_0 & (i_2_1_41_0 | (i_2_1_135_0 & i_2_1_136_0))))))) | (i_2_1_34_0 & ((~i_2_1_49_0 & (((i_2_1_136_0 | (~i_2_1_46_0 & i_2_1_135_0)) & (i_2_1_13_0 | (~i_2_1_54_0 & i_2_1_70_0))) | (i_2_1_41_0 & ~i_2_1_46_0 & (~i_2_1_54_0 | (i_2_1_70_0 & i_2_1_136_0))))) | (~i_2_1_54_0 & ((i_2_1_13_0 & ((i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_46_0 & i_2_1_70_0))) | (i_2_1_70_0 & i_2_1_135_0 & (i_2_1_136_0 | (i_2_1_41_0 & i_2_1_49_0))))))) | (i_2_1_13_0 & i_2_1_70_0 & ((~i_2_1_49_0 & i_2_1_135_0 & (~i_2_1_54_0 | (i_2_1_41_0 & ~i_2_1_46_0 & i_2_1_136_0))) | (~i_2_1_54_0 & i_2_1_136_0))))) | (~i_2_1_54_0 & ((~i_2_1_57_0 & ((i_2_1_32_0 & ((~i_2_1_38_0 & ((i_2_1_41_0 & i_2_1_70_0) | (i_2_1_13_0 & ~i_2_1_46_0 & i_2_1_51_0 & ~i_2_1_135_0))) | (i_2_1_136_0 & ((i_2_1_34_0 & (i_2_1_68_0 | (~i_2_1_41_0 & i_2_1_51_0 & i_2_1_135_0))) | (i_2_1_68_0 & ((~i_2_1_46_0 & i_2_1_135_0) | (~i_2_1_49_0 & (i_2_1_38_0 | (i_2_1_41_0 & i_2_1_135_0))))) | (~i_2_1_41_0 & i_2_1_49_0 & i_2_1_51_0 & i_2_1_70_0 & ~i_2_1_135_0))) | (i_2_1_38_0 & (((~i_2_1_46_0 | i_2_1_68_0) & (i_2_1_34_0 | i_2_1_41_0 | (~i_2_1_49_0 & i_2_1_70_0))) | (i_2_1_68_0 & (~i_2_1_46_0 | i_2_1_135_0)) | (i_2_1_13_0 & i_2_1_46_0))) | (i_2_1_41_0 & ((i_2_1_34_0 & i_2_1_68_0) | (i_2_1_13_0 & ~i_2_1_49_0))) | (i_2_1_68_0 & ((i_2_1_13_0 & (i_2_1_34_0 | i_2_1_135_0)) | (i_2_1_34_0 & ~i_2_1_46_0))) | (i_2_1_34_0 & i_2_1_135_0 & (~i_2_1_49_0 | i_2_1_70_0)))) | (((~i_2_1_46_0 & i_2_1_70_0) | (i_2_1_34_0 & i_2_1_41_0)) & ((i_2_1_38_0 & i_2_1_68_0) | (~i_2_1_49_0 & ~i_2_1_135_0 & i_2_1_136_0))) | (((i_2_1_34_0 & i_2_1_135_0) | (i_2_1_13_0 & i_2_1_38_0)) & ((~i_2_1_46_0 & i_2_1_68_0) | (i_2_1_41_0 & ~i_2_1_136_0))) | (i_2_1_68_0 & ((i_2_1_34_0 & ((i_2_1_41_0 & (i_2_1_70_0 | i_2_1_135_0)) | (i_2_1_135_0 & (i_2_1_13_0 | (~i_2_1_49_0 & i_2_1_136_0))) | ((i_2_1_38_0 | ~i_2_1_46_0 | ~i_2_1_49_0) & (i_2_1_13_0 | i_2_1_70_0)) | (~i_2_1_46_0 & (i_2_1_38_0 | ~i_2_1_49_0)) | (i_2_1_38_0 & (~i_2_1_49_0 | i_2_1_136_0)))) | (~i_2_1_46_0 & ((i_2_1_38_0 & (i_2_1_41_0 | (~i_2_1_49_0 & i_2_1_135_0))) | (~i_2_1_49_0 & ((i_2_1_135_0 & i_2_1_136_0) | (i_2_1_41_0 & i_2_1_70_0))) | (i_2_1_13_0 & (i_2_1_70_0 | i_2_1_135_0 | i_2_1_136_0)))) | (~i_2_1_49_0 & ((i_2_1_70_0 & ((i_2_1_38_0 & i_2_1_41_0) | (i_2_1_135_0 & ~i_2_1_136_0))) | (i_2_1_13_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_41_0 & ((i_2_1_70_0 & i_2_1_135_0) | ((i_2_1_135_0 | i_2_1_136_0) & (i_2_1_13_0 | i_2_1_38_0)))) | (i_2_1_38_0 & i_2_1_135_0 & (i_2_1_13_0 | i_2_1_136_0)))) | (i_2_1_38_0 & ((~i_2_1_49_0 & ((i_2_1_41_0 & (i_2_1_34_0 | (~i_2_1_46_0 & i_2_1_70_0))) | (i_2_1_70_0 & (i_2_1_135_0 | (~i_2_1_46_0 & i_2_1_136_0))))) | (~i_2_1_46_0 & ((~i_2_1_41_0 & i_2_1_135_0 & i_2_1_136_0) | (i_2_1_34_0 & (i_2_1_13_0 | i_2_1_70_0)))) | (i_2_1_13_0 & (i_2_1_70_0 | (~i_2_1_135_0 & i_2_1_136_0))))) | (~i_2_1_46_0 & ((~i_2_1_49_0 & ~i_2_1_70_0 & i_2_1_13_0 & ~i_2_1_34_0) | (i_2_1_34_0 & i_2_1_41_0 & i_2_1_136_0))) | (i_2_1_70_0 & ((i_2_1_13_0 & (i_2_1_34_0 | i_2_1_41_0)) | (i_2_1_136_0 & ((i_2_1_34_0 & i_2_1_135_0) | (i_2_1_41_0 & ~i_2_1_49_0))))) | (i_2_1_13_0 & i_2_1_34_0 & i_2_1_136_0))) | (i_2_1_32_0 & ((i_2_1_13_0 & ((~i_2_1_41_0 & ((i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_46_0 & ~i_2_1_49_0 & i_2_1_51_0 & ~i_2_1_70_0))) | (~i_2_1_49_0 & (i_2_1_136_0 | (i_2_1_34_0 & i_2_1_68_0))) | (i_2_1_135_0 & (i_2_1_70_0 | (i_2_1_41_0 & i_2_1_68_0))) | (i_2_1_41_0 & (i_2_1_38_0 | i_2_1_70_0)) | (i_2_1_38_0 & (i_2_1_70_0 | (i_2_1_34_0 & i_2_1_68_0))) | (i_2_1_34_0 & ((~i_2_1_46_0 & i_2_1_68_0) | (i_2_1_51_0 & i_2_1_70_0))) | (i_2_1_49_0 & i_2_1_68_0 & i_2_1_70_0))) | (i_2_1_135_0 & ((i_2_1_46_0 & ((i_2_1_70_0 & i_2_1_136_0) | (i_2_1_38_0 & i_2_1_41_0 & ~i_2_1_49_0 & ~i_2_1_70_0))) | (i_2_1_34_0 & ((i_2_1_38_0 & (i_2_1_41_0 | i_2_1_68_0)) | (i_2_1_41_0 & (i_2_1_70_0 | ((~i_2_1_49_0 | i_2_1_136_0) & (~i_2_1_46_0 | i_2_1_68_0)))) | (~i_2_1_49_0 & ((i_2_1_68_0 & i_2_1_136_0) | (i_2_1_51_0 & i_2_1_70_0))) | (i_2_1_70_0 & i_2_1_136_0) | (~i_2_1_46_0 & i_2_1_68_0))) | (i_2_1_38_0 & ((i_2_1_68_0 & i_2_1_136_0) | (~i_2_1_46_0 & i_2_1_70_0))) | (i_2_1_68_0 & ((i_2_1_70_0 & i_2_1_136_0) | (~i_2_1_49_0 & (i_2_1_70_0 | (~i_2_1_46_0 & i_2_1_136_0))))))) | (i_2_1_68_0 & ((i_2_1_41_0 & ((i_2_1_34_0 & (i_2_1_70_0 | (~i_2_1_49_0 & i_2_1_136_0))) | (~i_2_1_46_0 & (i_2_1_136_0 | (i_2_1_49_0 & i_2_1_51_0 & i_2_1_57_0))) | (i_2_1_38_0 & (i_2_1_49_0 | i_2_1_70_0 | i_2_1_136_0)))) | (i_2_1_136_0 & ((~i_2_1_49_0 & i_2_1_70_0) | (i_2_1_34_0 & i_2_1_38_0))) | (i_2_1_34_0 & ((~i_2_1_46_0 & ~i_2_1_49_0) | ((i_2_1_38_0 | i_2_1_70_0) & (~i_2_1_46_0 | ~i_2_1_49_0)))) | (i_2_1_38_0 & ~i_2_1_46_0 & ~i_2_1_49_0))) | (~i_2_1_46_0 & ((i_2_1_70_0 & ((i_2_1_34_0 & (i_2_1_38_0 | (i_2_1_41_0 & ~i_2_1_49_0))) | (i_2_1_38_0 & ~i_2_1_49_0 & i_2_1_136_0))) | (i_2_1_34_0 & ~i_2_1_49_0 & i_2_1_136_0))) | (i_2_1_70_0 & i_2_1_136_0 & i_2_1_41_0 & ~i_2_1_49_0))) | (i_2_1_38_0 & ((i_2_1_49_0 & ((i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_46_0 & i_2_1_70_0) | (i_2_1_13_0 & i_2_1_41_0 & i_2_1_51_0 & ~i_2_1_136_0))) | (i_2_1_13_0 & ((~i_2_1_49_0 & ((i_2_1_34_0 & i_2_1_68_0) | (~i_2_1_46_0 & ~i_2_1_70_0))) | (i_2_1_70_0 & (i_2_1_68_0 | (i_2_1_34_0 & ~i_2_1_46_0))) | (i_2_1_68_0 & ((i_2_1_34_0 & (~i_2_1_46_0 | i_2_1_135_0)) | (i_2_1_135_0 & (~i_2_1_46_0 | i_2_1_136_0)))) | (i_2_1_41_0 & i_2_1_135_0 & ~i_2_1_136_0))) | ((i_2_1_34_0 | ~i_2_1_46_0) & ((i_2_1_41_0 & i_2_1_70_0 & (i_2_1_68_0 | i_2_1_135_0)) | (i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_49_0 & i_2_1_68_0))) | (~i_2_1_46_0 & ((i_2_1_34_0 & (((i_2_1_68_0 | i_2_1_70_0) & (i_2_1_41_0 | ~i_2_1_49_0)) | (i_2_1_135_0 & (i_2_1_68_0 | (i_2_1_41_0 & i_2_1_136_0))) | (i_2_1_68_0 & (i_2_1_70_0 | i_2_1_136_0)))) | (i_2_1_41_0 & i_2_1_136_0 & (i_2_1_68_0 | i_2_1_70_0)) | (~i_2_1_49_0 & i_2_1_68_0 & i_2_1_70_0))) | (i_2_1_34_0 & ((i_2_1_68_0 & ((i_2_1_70_0 & i_2_1_135_0) | (i_2_1_41_0 & (~i_2_1_49_0 | (i_2_1_135_0 & i_2_1_136_0))))) | (~i_2_1_49_0 & i_2_1_70_0 & ~i_2_1_135_0))) | (i_2_1_68_0 & i_2_1_70_0 & (i_2_1_136_0 | (i_2_1_41_0 & i_2_1_135_0))))) | (i_2_1_34_0 & (((~i_2_1_49_0 | i_2_1_136_0) & ((i_2_1_41_0 & ((~i_2_1_46_0 & (i_2_1_68_0 | (i_2_1_70_0 & i_2_1_135_0))) | (i_2_1_68_0 & (i_2_1_13_0 | (i_2_1_70_0 & i_2_1_135_0))))) | (~i_2_1_46_0 & i_2_1_68_0 & i_2_1_70_0))) | (((~i_2_1_46_0 & (i_2_1_68_0 | (~i_2_1_49_0 & i_2_1_136_0))) | (~i_2_1_49_0 & i_2_1_68_0 & i_2_1_136_0)) & ((i_2_1_70_0 & i_2_1_135_0) | (i_2_1_41_0 & (i_2_1_70_0 | i_2_1_135_0)))) | (i_2_1_68_0 & ((~i_2_1_49_0 & ((i_2_1_13_0 & ~i_2_1_46_0) | ((i_2_1_135_0 | i_2_1_136_0) & (i_2_1_13_0 | ~i_2_1_46_0)))) | (i_2_1_13_0 & ~i_2_1_46_0 & (i_2_1_70_0 | i_2_1_135_0)))) | (i_2_1_13_0 & i_2_1_70_0 & (~i_2_1_49_0 | (~i_2_1_46_0 & i_2_1_135_0))))) | (i_2_1_70_0 & ((i_2_1_135_0 & ((i_2_1_13_0 & (i_2_1_41_0 | (~i_2_1_46_0 & i_2_1_68_0))) | (~i_2_1_46_0 & ~i_2_1_49_0 & i_2_1_68_0 & (i_2_1_41_0 | i_2_1_136_0)))) | (i_2_1_13_0 & ((~i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_49_0 & (i_2_1_136_0 | (~i_2_1_46_0 & i_2_1_68_0))))))) | (i_2_1_41_0 & i_2_1_136_0 & ((i_2_1_13_0 & ((~i_2_1_46_0 & i_2_1_51_0) | (~i_2_1_49_0 & i_2_1_68_0 & i_2_1_135_0))) | (i_2_1_68_0 & i_2_1_135_0 & ~i_2_1_46_0 & ~i_2_1_49_0))))) | (i_2_1_38_0 & ((~i_2_1_57_0 & ((i_2_1_136_0 & ((i_2_1_135_0 & ((i_2_1_32_0 & ((i_2_1_34_0 & (~i_2_1_46_0 | (~i_2_1_41_0 & ~i_2_1_70_0))) | (i_2_1_68_0 & (i_2_1_13_0 | (i_2_1_41_0 & ~i_2_1_49_0))) | (i_2_1_51_0 & ~i_2_1_70_0 & ~i_2_1_41_0 & ~i_2_1_46_0))) | (~i_2_1_49_0 & ((i_2_1_34_0 & i_2_1_68_0) | (i_2_1_41_0 & i_2_1_70_0))) | ((i_2_1_13_0 | i_2_1_34_0) & ((~i_2_1_46_0 & i_2_1_70_0) | (i_2_1_41_0 & i_2_1_68_0))) | (~i_2_1_46_0 & i_2_1_68_0 & (i_2_1_13_0 | i_2_1_41_0 | i_2_1_70_0)))) | (i_2_1_41_0 & ((~i_2_1_135_0 & ((i_2_1_13_0 & (~i_2_1_46_0 | ~i_2_1_49_0)) | (i_2_1_34_0 & i_2_1_70_0) | (~i_2_1_46_0 & ~i_2_1_49_0 & i_2_1_54_0))) | (i_2_1_68_0 & ((i_2_1_34_0 & ~i_2_1_49_0) | (~i_2_1_46_0 & i_2_1_70_0))))) | (i_2_1_70_0 & ((i_2_1_13_0 & (i_2_1_32_0 | ~i_2_1_49_0)) | (i_2_1_32_0 & (i_2_1_68_0 | (i_2_1_34_0 & ~i_2_1_46_0))) | (~i_2_1_46_0 & ~i_2_1_49_0 & i_2_1_68_0))) | (~i_2_1_49_0 & ((i_2_1_13_0 & (i_2_1_32_0 | ~i_2_1_46_0)) | (i_2_1_32_0 & ~i_2_1_46_0 & ~i_2_1_70_0))))) | (~i_2_1_49_0 & ((i_2_1_41_0 & ((i_2_1_32_0 & (i_2_1_34_0 | (i_2_1_54_0 & i_2_1_70_0))) | (i_2_1_34_0 & (i_2_1_70_0 | (i_2_1_135_0 & ~i_2_1_136_0))) | (i_2_1_68_0 & ((~i_2_1_46_0 & i_2_1_70_0) | (i_2_1_13_0 & i_2_1_135_0))) | (i_2_1_13_0 & (~i_2_1_46_0 | i_2_1_70_0)) | (~i_2_1_70_0 & i_2_1_135_0 & ~i_2_1_136_0 & ~i_2_1_46_0 & i_2_1_54_0))) | (i_2_1_68_0 & ((i_2_1_13_0 & (i_2_1_34_0 | (~i_2_1_46_0 & i_2_1_135_0))) | (~i_2_1_46_0 & (i_2_1_34_0 | (i_2_1_70_0 & (i_2_1_32_0 | i_2_1_135_0)))))) | (i_2_1_135_0 & ((i_2_1_32_0 & ~i_2_1_46_0 & ~i_2_1_70_0) | ((i_2_1_13_0 | i_2_1_34_0) & (i_2_1_32_0 | i_2_1_70_0)))) | (i_2_1_13_0 & i_2_1_32_0 & i_2_1_70_0))) | (i_2_1_70_0 & ((i_2_1_13_0 & (i_2_1_34_0 | (~i_2_1_46_0 & i_2_1_68_0))) | (i_2_1_135_0 & ((i_2_1_32_0 & ((i_2_1_41_0 & ~i_2_1_46_0) | (i_2_1_34_0 & ~i_2_1_136_0))) | (i_2_1_41_0 & i_2_1_49_0 & i_2_1_68_0 & ~i_2_1_136_0))) | (i_2_1_34_0 & i_2_1_68_0 & (i_2_1_32_0 | ~i_2_1_46_0)))) | (i_2_1_13_0 & ((i_2_1_41_0 & (i_2_1_34_0 | (i_2_1_32_0 & i_2_1_68_0))) | (i_2_1_68_0 & ((i_2_1_34_0 & ~i_2_1_46_0) | (i_2_1_32_0 & (i_2_1_34_0 | ~i_2_1_46_0)))))))) | (i_2_1_68_0 & ((i_2_1_70_0 & ((i_2_1_34_0 & ((i_2_1_13_0 & (~i_2_1_46_0 | ~i_2_1_49_0)) | (i_2_1_32_0 & (i_2_1_41_0 | (i_2_1_49_0 & ~i_2_1_135_0))) | (~i_2_1_46_0 & (i_2_1_41_0 | ~i_2_1_49_0 | i_2_1_135_0)) | (~i_2_1_41_0 & i_2_1_49_0 & i_2_1_57_0 & i_2_1_136_0))) | (i_2_1_32_0 & ((~i_2_1_49_0 & i_2_1_136_0) | (i_2_1_13_0 & ~i_2_1_46_0))) | (i_2_1_13_0 & ((~i_2_1_49_0 & (~i_2_1_46_0 | (i_2_1_41_0 & i_2_1_135_0))) | (i_2_1_41_0 & (~i_2_1_46_0 | i_2_1_136_0)) | (i_2_1_136_0 & (~i_2_1_46_0 | i_2_1_135_0)))) | (~i_2_1_46_0 & ((i_2_1_41_0 & ((i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_49_0 & (i_2_1_135_0 | i_2_1_136_0)))) | (~i_2_1_49_0 & i_2_1_135_0 & i_2_1_136_0))))) | (i_2_1_136_0 & ((i_2_1_32_0 & ((i_2_1_13_0 & (i_2_1_41_0 | ~i_2_1_46_0)) | (i_2_1_34_0 & (~i_2_1_46_0 | ~i_2_1_49_0)) | (~i_2_1_46_0 & ~i_2_1_49_0 & i_2_1_135_0))) | (i_2_1_135_0 & ((~i_2_1_46_0 & ((i_2_1_34_0 & i_2_1_41_0) | (i_2_1_13_0 & (i_2_1_41_0 | ~i_2_1_49_0)))) | (i_2_1_34_0 & i_2_1_41_0 & ~i_2_1_49_0))))) | (~i_2_1_46_0 & ~i_2_1_49_0 & ((i_2_1_13_0 & (i_2_1_34_0 | (i_2_1_41_0 & i_2_1_135_0))) | (i_2_1_34_0 & i_2_1_41_0) | (i_2_1_32_0 & (i_2_1_34_0 | i_2_1_41_0)))) | (i_2_1_32_0 & i_2_1_41_0 & i_2_1_51_0 & i_2_1_57_0 & i_2_1_135_0 & ~i_2_1_136_0))) | (~i_2_1_46_0 & ((i_2_1_13_0 & ((i_2_1_32_0 & ((i_2_1_135_0 & i_2_1_136_0) | (i_2_1_34_0 & i_2_1_51_0 & i_2_1_57_0))) | (i_2_1_41_0 & ~i_2_1_49_0 & ((~i_2_1_135_0 & i_2_1_136_0) | (i_2_1_70_0 & i_2_1_135_0))) | (~i_2_1_70_0 & i_2_1_135_0 & i_2_1_34_0 & i_2_1_57_0))) | (i_2_1_41_0 & ((i_2_1_32_0 & ((~i_2_1_49_0 & i_2_1_70_0) | (~i_2_1_70_0 & ~i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_34_0 & i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_34_0 & ~i_2_1_49_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_34_0 & ((~i_2_1_49_0 & ((i_2_1_32_0 & (i_2_1_13_0 | (i_2_1_57_0 & i_2_1_136_0))) | (i_2_1_136_0 & ((i_2_1_13_0 & (i_2_1_41_0 | i_2_1_135_0)) | (i_2_1_41_0 & i_2_1_70_0 & ~i_2_1_135_0))) | (i_2_1_135_0 & ~i_2_1_136_0 & i_2_1_41_0 & i_2_1_70_0))) | (i_2_1_13_0 & i_2_1_41_0 & (i_2_1_70_0 | i_2_1_135_0)))) | (i_2_1_32_0 & i_2_1_70_0 & ((i_2_1_13_0 & (i_2_1_41_0 | i_2_1_135_0)) | (~i_2_1_49_0 & i_2_1_135_0 & i_2_1_136_0))))) | (i_2_1_13_0 & ((i_2_1_32_0 & ((i_2_1_136_0 & ((i_2_1_49_0 & ((i_2_1_41_0 & i_2_1_70_0) | (i_2_1_34_0 & i_2_1_57_0 & i_2_1_68_0))) | (~i_2_1_49_0 & ((i_2_1_34_0 & (i_2_1_41_0 | ~i_2_1_57_0)) | (i_2_1_41_0 & ((~i_2_1_46_0 & i_2_1_57_0) | (~i_2_1_57_0 & i_2_1_68_0 & i_2_1_135_0))) | (i_2_1_70_0 & (~i_2_1_46_0 | i_2_1_68_0)) | (~i_2_1_46_0 & i_2_1_68_0 & (~i_2_1_57_0 | i_2_1_135_0)))) | (i_2_1_68_0 & ((i_2_1_41_0 & (i_2_1_70_0 | (~i_2_1_46_0 & ~i_2_1_57_0))) | (i_2_1_135_0 & (i_2_1_34_0 | (~i_2_1_46_0 & (~i_2_1_57_0 | i_2_1_70_0)))))))) | (i_2_1_34_0 & ((~i_2_1_46_0 & i_2_1_68_0 & (~i_2_1_49_0 | ~i_2_1_57_0)) | (~i_2_1_57_0 & (i_2_1_41_0 | (~i_2_1_49_0 & i_2_1_135_0))) | (~i_2_1_49_0 & (i_2_1_70_0 | (i_2_1_41_0 & ~i_2_1_68_0))) | (i_2_1_41_0 & ((i_2_1_135_0 & ~i_2_1_136_0) | (i_2_1_49_0 & i_2_1_51_0))))) | (i_2_1_70_0 & ((~i_2_1_57_0 & (i_2_1_41_0 | (~i_2_1_49_0 & i_2_1_135_0))) | (i_2_1_68_0 & ((i_2_1_41_0 & (i_2_1_135_0 | (~i_2_1_46_0 & ~i_2_1_49_0))) | (~i_2_1_46_0 & (~i_2_1_57_0 | (~i_2_1_49_0 & i_2_1_135_0))))))) | (~i_2_1_46_0 & ~i_2_1_49_0 & ~i_2_1_57_0 & i_2_1_68_0 & i_2_1_135_0))) | (i_2_1_70_0 & ((i_2_1_41_0 & ((i_2_1_135_0 & ((~i_2_1_46_0 & i_2_1_68_0 & (~i_2_1_49_0 | i_2_1_136_0)) | (~i_2_1_136_0 & (~i_2_1_57_0 | (i_2_1_34_0 & ~i_2_1_49_0))))) | (i_2_1_34_0 & i_2_1_68_0 & i_2_1_136_0) | ((i_2_1_34_0 | (~i_2_1_49_0 & i_2_1_136_0)) & (~i_2_1_57_0 | (~i_2_1_46_0 & i_2_1_68_0))))) | (~i_2_1_57_0 & ((i_2_1_34_0 & i_2_1_49_0 & i_2_1_68_0) | (~i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_46_0 & ~i_2_1_49_0))) | (i_2_1_68_0 & ((~i_2_1_46_0 & ((~i_2_1_49_0 & (i_2_1_34_0 | (i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_34_0 & (i_2_1_135_0 | i_2_1_136_0)))) | (i_2_1_34_0 & i_2_1_135_0 & i_2_1_136_0))))) | (i_2_1_135_0 & ((i_2_1_34_0 & ((i_2_1_41_0 & (~i_2_1_57_0 | (~i_2_1_49_0 & i_2_1_68_0 & i_2_1_136_0))) | (~i_2_1_46_0 & ((~i_2_1_49_0 & i_2_1_136_0) | (~i_2_1_57_0 & i_2_1_68_0))) | (~i_2_1_49_0 & ~i_2_1_57_0 & i_2_1_136_0))) | (~i_2_1_46_0 & i_2_1_68_0 & i_2_1_136_0 & ((~i_2_1_49_0 & ~i_2_1_57_0) | (i_2_1_41_0 & (~i_2_1_49_0 | ~i_2_1_57_0)))))) | (~i_2_1_49_0 & ~i_2_1_57_0 & i_2_1_68_0 & i_2_1_34_0 & ~i_2_1_46_0))) | (i_2_1_34_0 & ((i_2_1_41_0 & ((i_2_1_136_0 & ((i_2_1_32_0 & ((~i_2_1_46_0 & (~i_2_1_49_0 | (i_2_1_51_0 & i_2_1_70_0 & ~i_2_1_135_0))) | (~i_2_1_57_0 & ((~i_2_1_49_0 & i_2_1_68_0) | (i_2_1_51_0 & ~i_2_1_135_0))))) | (~i_2_1_46_0 & ((~i_2_1_57_0 & i_2_1_70_0) | (i_2_1_68_0 & ((i_2_1_70_0 & i_2_1_135_0) | (~i_2_1_49_0 & (i_2_1_70_0 | i_2_1_135_0)))))))) | (i_2_1_70_0 & ((i_2_1_32_0 & (~i_2_1_57_0 | (~i_2_1_46_0 & i_2_1_68_0))) | (i_2_1_135_0 & ((~i_2_1_57_0 & ~i_2_1_136_0) | (~i_2_1_46_0 & ~i_2_1_49_0 & i_2_1_68_0))))) | (~i_2_1_32_0 & ~i_2_1_46_0 & i_2_1_49_0 & ~i_2_1_57_0 & i_2_1_68_0 & ~i_2_1_135_0))) | (i_2_1_70_0 & ((~i_2_1_49_0 & ((i_2_1_68_0 & (((~i_2_1_46_0 | i_2_1_135_0) & (i_2_1_32_0 | ~i_2_1_57_0)) | (i_2_1_136_0 & (i_2_1_32_0 | (~i_2_1_46_0 & i_2_1_135_0))))) | (~i_2_1_57_0 & (i_2_1_136_0 | (i_2_1_32_0 & ~i_2_1_46_0))))) | (i_2_1_135_0 & i_2_1_136_0 & i_2_1_32_0 & i_2_1_68_0))) | (i_2_1_32_0 & ~i_2_1_46_0 & ~i_2_1_49_0 & ~i_2_1_57_0 & i_2_1_135_0))) | (~i_2_1_46_0 & ((i_2_1_68_0 & ((i_2_1_32_0 & ((~i_2_1_49_0 & ((~i_2_1_57_0 & ((i_2_1_70_0 & (i_2_1_135_0 | i_2_1_136_0)) | (i_2_1_41_0 & (i_2_1_70_0 | (i_2_1_135_0 & i_2_1_136_0))))) | (i_2_1_41_0 & i_2_1_70_0 & i_2_1_135_0))) | (i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0 & (i_2_1_41_0 | ~i_2_1_57_0)))) | (i_2_1_41_0 & ~i_2_1_49_0 & ~i_2_1_57_0 & i_2_1_70_0 & (i_2_1_135_0 | i_2_1_136_0)))) | (i_2_1_32_0 & i_2_1_41_0 & ~i_2_1_49_0 & ~i_2_1_57_0 & i_2_1_70_0 & i_2_1_135_0))) | (~i_2_1_49_0 & ~i_2_1_57_0 & i_2_1_32_0 & i_2_1_41_0 & i_2_1_135_0 & i_2_1_136_0 & i_2_1_68_0 & i_2_1_70_0))) | (~i_2_1_54_0 & ((~i_2_1_49_0 & ((i_2_1_32_0 & ((~i_2_1_38_0 & ((i_2_1_13_0 & ~i_2_1_46_0 & ~i_2_1_70_0 & i_2_1_135_0) | (i_2_1_34_0 & i_2_1_41_0 & ~i_2_1_51_0 & ~i_2_1_57_0 & ~i_2_1_136_0))) | (~i_2_1_57_0 & ((~i_2_1_51_0 & ((~i_2_1_41_0 & ((i_2_1_13_0 & i_2_1_135_0 & i_2_1_136_0) | (i_2_1_68_0 & i_2_1_70_0 & ~i_2_1_136_0))) | ((i_2_1_34_0 | (i_2_1_41_0 & i_2_1_136_0)) & ((i_2_1_70_0 & ~i_2_1_135_0) | (i_2_1_68_0 & (i_2_1_38_0 | i_2_1_135_0)))) | (i_2_1_136_0 & ((i_2_1_34_0 & (i_2_1_70_0 | (i_2_1_38_0 & i_2_1_41_0))) | (~i_2_1_46_0 & (i_2_1_41_0 | i_2_1_135_0 | (i_2_1_38_0 & i_2_1_70_0))))) | (i_2_1_34_0 & ((i_2_1_13_0 & i_2_1_68_0) | (i_2_1_41_0 & i_2_1_135_0))) | (i_2_1_13_0 & i_2_1_68_0 & (i_2_1_38_0 | i_2_1_41_0)))) | (i_2_1_136_0 & ((i_2_1_51_0 & ((i_2_1_13_0 & i_2_1_41_0) | (~i_2_1_46_0 & i_2_1_68_0 & ~i_2_1_135_0))) | (i_2_1_13_0 & (i_2_1_34_0 | (i_2_1_38_0 & i_2_1_68_0))) | (i_2_1_38_0 & (((i_2_1_34_0 | i_2_1_70_0) & (i_2_1_68_0 | (i_2_1_41_0 & i_2_1_135_0))) | (i_2_1_41_0 & i_2_1_68_0 & i_2_1_135_0))) | (i_2_1_135_0 & ((~i_2_1_46_0 & i_2_1_70_0) | (i_2_1_41_0 & (~i_2_1_46_0 | (i_2_1_68_0 & i_2_1_70_0))))))) | (i_2_1_68_0 & ((i_2_1_70_0 & (~i_2_1_46_0 | (i_2_1_38_0 & i_2_1_41_0))) | (~i_2_1_46_0 & (i_2_1_41_0 | (i_2_1_135_0 & ~i_2_1_136_0))) | (i_2_1_38_0 & (i_2_1_13_0 | i_2_1_34_0) & (i_2_1_41_0 | i_2_1_135_0)) | (i_2_1_13_0 & i_2_1_34_0 & i_2_1_135_0))) | (i_2_1_70_0 & (((i_2_1_41_0 | ~i_2_1_46_0) & (i_2_1_13_0 | (i_2_1_34_0 & i_2_1_38_0))) | (i_2_1_41_0 & ~i_2_1_46_0) | (i_2_1_34_0 & i_2_1_51_0 & i_2_1_135_0))) | (i_2_1_13_0 & i_2_1_34_0 & i_2_1_41_0))) | (i_2_1_68_0 & ((i_2_1_70_0 & ((i_2_1_51_0 & ((i_2_1_38_0 & i_2_1_136_0) | (i_2_1_135_0 & ~i_2_1_136_0 & i_2_1_41_0 & i_2_1_57_0))) | (i_2_1_34_0 & ((i_2_1_38_0 & (~i_2_1_51_0 | i_2_1_135_0)) | i_2_1_13_0 | ~i_2_1_46_0 | (~i_2_1_51_0 & (i_2_1_41_0 | i_2_1_135_0)))) | (i_2_1_41_0 & ~i_2_1_51_0 & i_2_1_136_0))) | (~i_2_1_51_0 & ((~i_2_1_46_0 & (i_2_1_41_0 | (i_2_1_34_0 & i_2_1_135_0))) | (i_2_1_41_0 & ((i_2_1_13_0 & (i_2_1_34_0 | i_2_1_136_0)) | (i_2_1_38_0 & i_2_1_135_0 & i_2_1_136_0) | (i_2_1_34_0 & (i_2_1_38_0 | i_2_1_136_0)))) | (i_2_1_135_0 & ((i_2_1_34_0 & i_2_1_38_0) | (i_2_1_13_0 & (i_2_1_34_0 | i_2_1_38_0)))))) | (i_2_1_34_0 & ((i_2_1_13_0 & i_2_1_38_0) | ((i_2_1_13_0 | i_2_1_38_0) & (~i_2_1_46_0 | (i_2_1_135_0 & (i_2_1_41_0 | i_2_1_136_0)))))) | (i_2_1_13_0 & i_2_1_41_0 & ((~i_2_1_135_0 & i_2_1_136_0) | (i_2_1_38_0 & i_2_1_135_0))))) | (i_2_1_13_0 & ((~i_2_1_46_0 & ((i_2_1_34_0 & i_2_1_135_0) | (~i_2_1_51_0 & i_2_1_70_0 & ~i_2_1_135_0))) | (i_2_1_34_0 & ((i_2_1_41_0 & ~i_2_1_51_0 & i_2_1_136_0) | (i_2_1_38_0 & i_2_1_135_0))) | (i_2_1_38_0 & ((i_2_1_41_0 & i_2_1_70_0) | (~i_2_1_51_0 & i_2_1_57_0 & i_2_1_136_0))) | (i_2_1_70_0 & i_2_1_135_0 & (i_2_1_41_0 | (~i_2_1_34_0 & i_2_1_46_0 & ~i_2_1_51_0 & i_2_1_57_0))))) | (i_2_1_34_0 & ((i_2_1_41_0 & ((i_2_1_136_0 & ((i_2_1_38_0 & (i_2_1_70_0 | (~i_2_1_51_0 & i_2_1_135_0))) | ~i_2_1_46_0 | (~i_2_1_51_0 & i_2_1_70_0 & i_2_1_135_0))) | (~i_2_1_46_0 & i_2_1_70_0 & i_2_1_135_0))) | (~i_2_1_46_0 & ((i_2_1_70_0 & i_2_1_136_0) | (i_2_1_38_0 & i_2_1_135_0))))) | (i_2_1_41_0 & ~i_2_1_46_0 & ~i_2_1_51_0 & i_2_1_70_0 & i_2_1_135_0))) | (i_2_1_135_0 & ((i_2_1_70_0 & ((~i_2_1_32_0 & i_2_1_47_0 & ((i_2_1_68_0 & i_2_1_136_0 & ~i_2_1_41_0 & ~i_2_1_57_0) | (i_2_1_13_0 & ~i_2_1_46_0 & i_2_1_51_0 & ~i_2_1_68_0 & ~i_2_1_136_0))) | (i_2_1_13_0 & ((i_2_1_38_0 & (~i_2_1_41_0 | i_2_1_68_0)) | (~i_2_1_57_0 & (i_2_1_34_0 | (i_2_1_51_0 & ~i_2_1_68_0))) | (i_2_1_34_0 & ((i_2_1_68_0 & (i_2_1_41_0 | ~i_2_1_51_0)) | (~i_2_1_41_0 & i_2_1_136_0))))) | (~i_2_1_51_0 & ((~i_2_1_46_0 & ((i_2_1_68_0 & ~i_2_1_136_0) | (i_2_1_136_0 & (i_2_1_38_0 | i_2_1_41_0)))) | (i_2_1_38_0 & (i_2_1_68_0 | (i_2_1_41_0 & ~i_2_1_57_0 & ~i_2_1_136_0))) | (~i_2_1_57_0 & (i_2_1_68_0 | (i_2_1_34_0 & i_2_1_41_0))))) | (i_2_1_34_0 & ((i_2_1_68_0 & ((i_2_1_38_0 & (i_2_1_41_0 | ~i_2_1_57_0)) | (i_2_1_136_0 & (i_2_1_41_0 | ~i_2_1_46_0)))) | (~i_2_1_57_0 & (~i_2_1_46_0 | (i_2_1_38_0 & i_2_1_136_0))))) | (i_2_1_38_0 & i_2_1_41_0 & ~i_2_1_46_0 & ~i_2_1_57_0 & i_2_1_136_0))) | (i_2_1_68_0 & (((~i_2_1_51_0 | i_2_1_136_0) & ((i_2_1_34_0 & ((i_2_1_38_0 & i_2_1_41_0) | (i_2_1_13_0 & (i_2_1_38_0 | i_2_1_41_0)))) | (~i_2_1_41_0 & ~i_2_1_57_0 & ~i_2_1_32_0 & i_2_1_38_0))) | (~i_2_1_46_0 & ((i_2_1_13_0 & (i_2_1_34_0 | i_2_1_136_0)) | (i_2_1_34_0 & (i_2_1_41_0 | (~i_2_1_51_0 & i_2_1_136_0))) | (i_2_1_38_0 & (i_2_1_41_0 | ~i_2_1_51_0)) | (i_2_1_41_0 & ~i_2_1_136_0 & (~i_2_1_51_0 | ~i_2_1_57_0)))) | (~i_2_1_51_0 & i_2_1_136_0 & ((i_2_1_38_0 & ~i_2_1_57_0) | (i_2_1_13_0 & i_2_1_34_0))) | (i_2_1_41_0 & ~i_2_1_57_0 & ((i_2_1_34_0 & i_2_1_38_0) | (i_2_1_13_0 & (i_2_1_34_0 | i_2_1_38_0)))))) | (i_2_1_34_0 & ((~i_2_1_57_0 & ((i_2_1_13_0 & ((i_2_1_38_0 & i_2_1_41_0) | (~i_2_1_41_0 & i_2_1_136_0))) | (i_2_1_38_0 & (~i_2_1_46_0 | (~i_2_1_51_0 & i_2_1_136_0))))) | (i_2_1_38_0 & ~i_2_1_46_0 & (i_2_1_41_0 | i_2_1_136_0)))) | (i_2_1_38_0 & i_2_1_41_0 & ~i_2_1_46_0 & ~i_2_1_51_0 & i_2_1_136_0))) | (~i_2_1_46_0 & ((i_2_1_136_0 & ((i_2_1_13_0 & ((i_2_1_47_0 & ~i_2_1_70_0) | (~i_2_1_51_0 & ~i_2_1_135_0))) | (i_2_1_38_0 & ((~i_2_1_57_0 & i_2_1_68_0) | (i_2_1_34_0 & ~i_2_1_70_0))) | (i_2_1_41_0 & ((~i_2_1_51_0 & ((i_2_1_68_0 & ~i_2_1_135_0) | (i_2_1_47_0 & i_2_1_70_0))) | (i_2_1_68_0 & ~i_2_1_135_0 & (~i_2_1_57_0 | i_2_1_70_0)))))) | (i_2_1_38_0 & ((i_2_1_41_0 & ((~i_2_1_57_0 & i_2_1_68_0 & i_2_1_70_0) | (i_2_1_34_0 & i_2_1_57_0 & ~i_2_1_70_0))) | (((~i_2_1_57_0 & i_2_1_68_0) | (i_2_1_34_0 & (i_2_1_68_0 | i_2_1_70_0))) & (i_2_1_13_0 | ~i_2_1_51_0)) | (i_2_1_68_0 & ((i_2_1_34_0 & (~i_2_1_57_0 | i_2_1_70_0)) | (i_2_1_13_0 & i_2_1_70_0))))) | (i_2_1_13_0 & ((~i_2_1_51_0 & (~i_2_1_57_0 | (i_2_1_34_0 & i_2_1_68_0))) | (i_2_1_68_0 & (i_2_1_41_0 | (i_2_1_34_0 & (~i_2_1_57_0 | i_2_1_70_0)))))) | (i_2_1_70_0 & ((i_2_1_41_0 & ((~i_2_1_51_0 & (i_2_1_68_0 | (i_2_1_34_0 & ~i_2_1_135_0))) | (i_2_1_34_0 & (~i_2_1_57_0 | i_2_1_68_0)))) | (i_2_1_34_0 & ~i_2_1_57_0 & i_2_1_68_0))))) | (i_2_1_34_0 & ((i_2_1_38_0 & ((i_2_1_41_0 & ((~i_2_1_51_0 & (i_2_1_13_0 | (~i_2_1_57_0 & i_2_1_68_0))) | (i_2_1_13_0 & (i_2_1_68_0 | (~i_2_1_57_0 & i_2_1_70_0))) | (~i_2_1_57_0 & i_2_1_68_0 & (i_2_1_70_0 | i_2_1_136_0)))) | (i_2_1_68_0 & ((~i_2_1_51_0 & i_2_1_136_0) | (i_2_1_13_0 & (~i_2_1_57_0 | i_2_1_70_0)))) | (~i_2_1_32_0 & ~i_2_1_41_0 & i_2_1_51_0 & ~i_2_1_57_0 & i_2_1_70_0 & i_2_1_136_0))) | (i_2_1_68_0 & i_2_1_136_0 & ((i_2_1_41_0 & ((i_2_1_13_0 & (~i_2_1_57_0 | i_2_1_70_0)) | (~i_2_1_51_0 & ~i_2_1_57_0))) | (~i_2_1_51_0 & ~i_2_1_57_0 & ~i_2_1_135_0))))) | (i_2_1_13_0 & ~i_2_1_51_0 & ((i_2_1_68_0 & i_2_1_70_0 & i_2_1_136_0) | (i_2_1_41_0 & ((~i_2_1_57_0 & i_2_1_68_0 & i_2_1_136_0) | (i_2_1_38_0 & (i_2_1_68_0 | (~i_2_1_57_0 & i_2_1_136_0))))))))) | (~i_2_1_57_0 & ((i_2_1_70_0 & ((~i_2_1_51_0 & ((i_2_1_13_0 & ((~i_2_1_32_0 & (i_2_1_34_0 | (i_2_1_135_0 & ~i_2_1_136_0))) | (i_2_1_41_0 & i_2_1_135_0 & (i_2_1_38_0 | (i_2_1_32_0 & i_2_1_136_0))) | (i_2_1_38_0 & (i_2_1_34_0 | ~i_2_1_46_0)) | (~i_2_1_34_0 & ~i_2_1_38_0 & ~i_2_1_41_0 & i_2_1_46_0 & ~i_2_1_135_0))) | (~i_2_1_46_0 & ((i_2_1_32_0 & ((i_2_1_135_0 & i_2_1_136_0) | (i_2_1_34_0 & i_2_1_38_0))) | (i_2_1_38_0 & ((i_2_1_41_0 & i_2_1_136_0) | (i_2_1_34_0 & (i_2_1_41_0 | i_2_1_136_0)))) | (i_2_1_68_0 & (i_2_1_135_0 | i_2_1_136_0)))) | (i_2_1_68_0 & ((i_2_1_38_0 & i_2_1_41_0) | (i_2_1_32_0 & ~i_2_1_38_0 & i_2_1_49_0))) | (i_2_1_32_0 & i_2_1_41_0 & ((i_2_1_38_0 & i_2_1_135_0 & i_2_1_136_0) | (i_2_1_34_0 & (i_2_1_38_0 | (i_2_1_135_0 & i_2_1_136_0))))) | (i_2_1_135_0 & i_2_1_136_0 & i_2_1_34_0 & i_2_1_38_0))) | (i_2_1_32_0 & ((~i_2_1_38_0 & ((~i_2_1_46_0 & i_2_1_68_0) | (i_2_1_34_0 & ~i_2_1_41_0 & i_2_1_46_0 & ~i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_34_0 & ((i_2_1_68_0 & (i_2_1_38_0 | i_2_1_41_0)) | (i_2_1_38_0 & (i_2_1_135_0 | i_2_1_136_0) & (i_2_1_41_0 | ~i_2_1_46_0)) | (i_2_1_41_0 & (i_2_1_13_0 | ~i_2_1_46_0)))) | (i_2_1_13_0 & ((i_2_1_38_0 & i_2_1_136_0) | (~i_2_1_41_0 & i_2_1_68_0))))) | (i_2_1_68_0 & ((i_2_1_38_0 & ((i_2_1_13_0 & (i_2_1_41_0 | ~i_2_1_46_0)) | (i_2_1_34_0 & ~i_2_1_46_0) | (i_2_1_135_0 & (i_2_1_136_0 | (~i_2_1_34_0 & i_2_1_49_0))))) | (i_2_1_13_0 & ((i_2_1_41_0 & i_2_1_136_0) | (i_2_1_34_0 & ~i_2_1_135_0))) | (i_2_1_41_0 & ((~i_2_1_46_0 & i_2_1_136_0) | (i_2_1_34_0 & (i_2_1_135_0 | i_2_1_136_0)))) | (~i_2_1_46_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_34_0 & i_2_1_38_0 & ((i_2_1_13_0 & (~i_2_1_46_0 | i_2_1_135_0)) | (~i_2_1_46_0 & ((i_2_1_135_0 & i_2_1_136_0) | (i_2_1_41_0 & (i_2_1_135_0 | i_2_1_136_0)))))))) | (i_2_1_68_0 & ((i_2_1_34_0 & ((~i_2_1_46_0 & ((i_2_1_13_0 & (i_2_1_32_0 | i_2_1_38_0)) | (~i_2_1_135_0 & (i_2_1_136_0 | (~i_2_1_32_0 & i_2_1_49_0 & ~i_2_1_51_0))) | i_2_1_41_0 | (i_2_1_38_0 & i_2_1_135_0))) | (i_2_1_13_0 & (((i_2_1_38_0 | (i_2_1_135_0 & i_2_1_136_0)) & (i_2_1_32_0 | i_2_1_41_0)) | (~i_2_1_51_0 & (i_2_1_38_0 | (i_2_1_32_0 & i_2_1_135_0))) | (i_2_1_38_0 & (i_2_1_135_0 | i_2_1_136_0)))) | (i_2_1_32_0 & ((i_2_1_41_0 & (i_2_1_135_0 | i_2_1_136_0)) | (i_2_1_38_0 & ((i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_51_0 & (i_2_1_41_0 | i_2_1_136_0)))))) | (i_2_1_135_0 & ((i_2_1_38_0 & i_2_1_136_0 & (i_2_1_41_0 | ~i_2_1_51_0)) | (i_2_1_41_0 & ~i_2_1_51_0 & ~i_2_1_136_0))))) | (i_2_1_135_0 & ((i_2_1_32_0 & ((i_2_1_41_0 & ((i_2_1_13_0 & ((i_2_1_51_0 & ~i_2_1_136_0) | (~i_2_1_51_0 & i_2_1_136_0))) | (i_2_1_38_0 & ~i_2_1_51_0))) | (~i_2_1_51_0 & ~i_2_1_136_0 & i_2_1_38_0 & i_2_1_49_0))) | (~i_2_1_46_0 & ((i_2_1_13_0 & ~i_2_1_51_0) | (i_2_1_41_0 & i_2_1_49_0 & i_2_1_136_0))))) | (i_2_1_38_0 & ((i_2_1_13_0 & ((i_2_1_41_0 & (~i_2_1_51_0 | i_2_1_136_0)) | (i_2_1_32_0 & ~i_2_1_46_0) | (~i_2_1_51_0 & i_2_1_136_0))) | (~i_2_1_46_0 & i_2_1_47_0 & i_2_1_136_0))))) | (i_2_1_32_0 & ((i_2_1_34_0 & ((i_2_1_136_0 & ((~i_2_1_51_0 & ((i_2_1_13_0 & (i_2_1_41_0 | ~i_2_1_135_0)) | ~i_2_1_46_0 | (i_2_1_38_0 & i_2_1_41_0 & i_2_1_135_0))) | (i_2_1_41_0 & ~i_2_1_46_0 & ~i_2_1_135_0))) | (~i_2_1_46_0 & ((i_2_1_13_0 & i_2_1_38_0) | (i_2_1_41_0 & i_2_1_135_0 & ~i_2_1_136_0))) | (i_2_1_13_0 & i_2_1_38_0 & ((~i_2_1_51_0 & i_2_1_135_0) | (i_2_1_41_0 & (~i_2_1_51_0 | i_2_1_135_0)))))) | (i_2_1_38_0 & i_2_1_41_0 & ~i_2_1_51_0 & i_2_1_135_0 & (~i_2_1_46_0 | (i_2_1_13_0 & i_2_1_136_0))))) | (i_2_1_38_0 & i_2_1_135_0 & ((i_2_1_13_0 & (~i_2_1_46_0 | (i_2_1_34_0 & i_2_1_41_0 & ~i_2_1_51_0))) | (~i_2_1_46_0 & i_2_1_136_0 & i_2_1_34_0 & i_2_1_41_0))) | (i_2_1_13_0 & ~i_2_1_34_0 & i_2_1_41_0 & ~i_2_1_46_0))) | (i_2_1_13_0 & ((~i_2_1_46_0 & ((~i_2_1_32_0 & ((i_2_1_38_0 & i_2_1_57_0 & i_2_1_136_0) | (i_2_1_34_0 & i_2_1_41_0 & i_2_1_49_0 & i_2_1_70_0 & ~i_2_1_135_0 & ~i_2_1_136_0))) | (i_2_1_32_0 & ((i_2_1_41_0 & (i_2_1_135_0 | (~i_2_1_51_0 & i_2_1_70_0))) | (i_2_1_34_0 & ((i_2_1_38_0 & (i_2_1_68_0 | i_2_1_70_0)) | (~i_2_1_51_0 & (i_2_1_68_0 | (i_2_1_70_0 & i_2_1_135_0))))) | (~i_2_1_51_0 & ((i_2_1_38_0 & i_2_1_68_0) | (~i_2_1_34_0 & i_2_1_136_0))) | (i_2_1_135_0 & (i_2_1_136_0 | (i_2_1_51_0 & i_2_1_68_0))))) | (i_2_1_34_0 & ((i_2_1_136_0 & ((i_2_1_68_0 & ~i_2_1_135_0) | (i_2_1_41_0 & i_2_1_70_0 & i_2_1_135_0))) | (i_2_1_41_0 & (i_2_1_68_0 | (i_2_1_38_0 & i_2_1_57_0))) | (i_2_1_68_0 & ((i_2_1_38_0 & (i_2_1_70_0 | i_2_1_135_0)) | (i_2_1_135_0 & (~i_2_1_51_0 | i_2_1_70_0)))))) | (i_2_1_41_0 & i_2_1_68_0 & (i_2_1_70_0 | i_2_1_136_0)))) | (i_2_1_32_0 & ((i_2_1_38_0 & ((i_2_1_70_0 & ((i_2_1_34_0 & i_2_1_135_0) | (~i_2_1_51_0 & i_2_1_136_0))) | (i_2_1_34_0 & ((~i_2_1_51_0 & (i_2_1_68_0 | (i_2_1_41_0 & i_2_1_135_0))) | ((i_2_1_68_0 | i_2_1_136_0) & (i_2_1_41_0 | i_2_1_135_0)) | (i_2_1_51_0 & i_2_1_57_0 & i_2_1_136_0))) | (i_2_1_68_0 & i_2_1_135_0 & (i_2_1_136_0 | (i_2_1_41_0 & ~i_2_1_51_0))))) | (i_2_1_34_0 & ((i_2_1_68_0 & (((i_2_1_70_0 | (i_2_1_135_0 & i_2_1_136_0)) & (i_2_1_41_0 | ~i_2_1_51_0)) | (i_2_1_41_0 & ~i_2_1_51_0 & i_2_1_135_0))) | (i_2_1_70_0 & i_2_1_135_0 & i_2_1_41_0 & ~i_2_1_51_0))) | (i_2_1_68_0 & i_2_1_70_0 & i_2_1_41_0 & ~i_2_1_51_0))) | (i_2_1_34_0 & ((i_2_1_38_0 & ((i_2_1_70_0 & (i_2_1_136_0 | ((i_2_1_41_0 | i_2_1_135_0) & (~i_2_1_51_0 | i_2_1_68_0)))) | (i_2_1_41_0 & i_2_1_68_0 & (~i_2_1_51_0 | i_2_1_136_0)))) | (i_2_1_41_0 & i_2_1_68_0 & ((i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_51_0 & (i_2_1_70_0 | i_2_1_136_0)))))) | (i_2_1_68_0 & i_2_1_70_0 & i_2_1_38_0 & ~i_2_1_51_0))) | (~i_2_1_46_0 & ((i_2_1_68_0 & ((i_2_1_136_0 & ((i_2_1_38_0 & (~i_2_1_51_0 | (i_2_1_34_0 & i_2_1_135_0))) | (i_2_1_70_0 & ((i_2_1_41_0 & ((~i_2_1_51_0 & ~i_2_1_135_0) | (i_2_1_49_0 & i_2_1_51_0 & i_2_1_135_0))) | (~i_2_1_51_0 & (i_2_1_32_0 | i_2_1_34_0)))) | (i_2_1_32_0 & i_2_1_34_0 & (i_2_1_135_0 | (i_2_1_49_0 & i_2_1_51_0))))) | (i_2_1_70_0 & ((i_2_1_34_0 & ((i_2_1_38_0 & i_2_1_41_0) | (i_2_1_32_0 & ~i_2_1_51_0))) | (i_2_1_38_0 & ((~i_2_1_51_0 & i_2_1_57_0) | (i_2_1_49_0 & (i_2_1_135_0 | (i_2_1_32_0 & i_2_1_57_0))))) | (i_2_1_32_0 & (i_2_1_41_0 | (i_2_1_47_0 & i_2_1_49_0 & i_2_1_135_0))))) | (i_2_1_32_0 & i_2_1_135_0 & ((i_2_1_41_0 & ~i_2_1_136_0) | (i_2_1_38_0 & i_2_1_49_0))))) | (i_2_1_38_0 & ((i_2_1_32_0 & ((i_2_1_34_0 & i_2_1_135_0 & i_2_1_136_0) | (i_2_1_70_0 & ((~i_2_1_51_0 & ((i_2_1_34_0 & i_2_1_136_0) | (i_2_1_49_0 & (i_2_1_135_0 | (i_2_1_41_0 & i_2_1_57_0))))) | (i_2_1_41_0 & ((i_2_1_135_0 & i_2_1_136_0) | (i_2_1_34_0 & (i_2_1_135_0 | i_2_1_136_0)))))))) | (i_2_1_41_0 & ((i_2_1_34_0 & i_2_1_136_0 & (~i_2_1_51_0 | (i_2_1_70_0 & i_2_1_135_0))) | (i_2_1_135_0 & ~i_2_1_136_0 & ~i_2_1_32_0 & ~i_2_1_51_0))))) | (~i_2_1_51_0 & i_2_1_70_0 & i_2_1_135_0 & i_2_1_32_0 & i_2_1_34_0 & i_2_1_41_0))) | (i_2_1_41_0 & ((i_2_1_70_0 & ((i_2_1_34_0 & ((i_2_1_32_0 & ((i_2_1_68_0 & i_2_1_136_0) | (i_2_1_38_0 & (i_2_1_68_0 | (~i_2_1_51_0 & i_2_1_135_0 & i_2_1_136_0))))) | (~i_2_1_51_0 & i_2_1_68_0 & (i_2_1_135_0 | i_2_1_136_0)))) | (i_2_1_38_0 & i_2_1_68_0 & ((~i_2_1_135_0 & i_2_1_136_0) | (i_2_1_32_0 & ~i_2_1_51_0))))) | (i_2_1_34_0 & i_2_1_38_0 & ~i_2_1_51_0 & i_2_1_68_0 & i_2_1_136_0))) | (i_2_1_68_0 & i_2_1_70_0 & i_2_1_136_0 & i_2_1_32_0 & i_2_1_34_0 & ~i_2_1_51_0))) | (i_2_1_13_0 & ((i_2_1_38_0 & ((i_2_1_32_0 & ((~i_2_1_46_0 & ((i_2_1_34_0 & (i_2_1_135_0 | (~i_2_1_51_0 & i_2_1_70_0))) | (i_2_1_41_0 & (~i_2_1_49_0 | (~i_2_1_51_0 & i_2_1_70_0 & i_2_1_136_0))) | (~i_2_1_70_0 & ((i_2_1_47_0 & ((i_2_1_57_0 & i_2_1_68_0 & ~i_2_1_49_0 & i_2_1_51_0) | (~i_2_1_41_0 & i_2_1_49_0 & ~i_2_1_51_0 & ~i_2_1_68_0 & i_2_1_136_0))) | (~i_2_1_49_0 & i_2_1_54_0 & i_2_1_57_0 & i_2_1_135_0))) | (~i_2_1_51_0 & ((~i_2_1_57_0 & i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_49_0 & i_2_1_68_0 & i_2_1_70_0))) | (i_2_1_68_0 & i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_49_0 & ((i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0) | (i_2_1_68_0 & (i_2_1_136_0 | (~i_2_1_57_0 & i_2_1_70_0))))))) | (i_2_1_34_0 & ((~i_2_1_49_0 & ((i_2_1_70_0 & (~i_2_1_57_0 | (i_2_1_41_0 & i_2_1_51_0 & ~i_2_1_135_0))) | (i_2_1_51_0 & ((~i_2_1_57_0 & i_2_1_135_0) | (~i_2_1_41_0 & i_2_1_136_0))) | (~i_2_1_51_0 & ((i_2_1_41_0 & i_2_1_68_0) | (~i_2_1_41_0 & ((~i_2_1_57_0 & ~i_2_1_135_0 & ~i_2_1_136_0) | (i_2_1_57_0 & i_2_1_135_0))))) | (i_2_1_135_0 & i_2_1_136_0) | (i_2_1_41_0 & i_2_1_68_0 & (~i_2_1_57_0 | i_2_1_135_0)))) | (~i_2_1_57_0 & ((~i_2_1_51_0 & i_2_1_70_0 & i_2_1_136_0) | (i_2_1_135_0 & ((i_2_1_41_0 & (i_2_1_68_0 | (~i_2_1_51_0 & i_2_1_136_0))) | (i_2_1_70_0 & i_2_1_136_0) | (i_2_1_68_0 & (~i_2_1_51_0 | i_2_1_136_0)))))) | (i_2_1_68_0 & ((i_2_1_49_0 & i_2_1_70_0) | (~i_2_1_51_0 & i_2_1_135_0 & i_2_1_136_0))))) | (~i_2_1_49_0 & ((i_2_1_41_0 & ((~i_2_1_51_0 & ((i_2_1_68_0 & (i_2_1_70_0 | (i_2_1_135_0 & i_2_1_136_0))) | (~i_2_1_57_0 & ((i_2_1_70_0 & i_2_1_136_0) | (i_2_1_68_0 & i_2_1_135_0))))) | (i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_57_0 & i_2_1_68_0))) | (i_2_1_68_0 & i_2_1_136_0 & ((i_2_1_51_0 & i_2_1_70_0) | (~i_2_1_51_0 & ~i_2_1_57_0 & i_2_1_135_0))))) | (~i_2_1_57_0 & i_2_1_68_0 & ((~i_2_1_51_0 & i_2_1_70_0 & ~i_2_1_135_0) | (i_2_1_41_0 & (i_2_1_70_0 | (~i_2_1_51_0 & i_2_1_135_0 & i_2_1_136_0))))))) | (~i_2_1_49_0 & ((i_2_1_70_0 & ((~i_2_1_41_0 & ((i_2_1_34_0 & ~i_2_1_51_0) | (~i_2_1_46_0 & ~i_2_1_57_0 & i_2_1_135_0))) | (i_2_1_41_0 & ((~i_2_1_46_0 & ~i_2_1_51_0 & i_2_1_136_0) | (i_2_1_68_0 & ((i_2_1_34_0 & (~i_2_1_57_0 | i_2_1_135_0)) | (~i_2_1_46_0 & (i_2_1_135_0 | i_2_1_136_0)) | (i_2_1_136_0 & (~i_2_1_51_0 | (~i_2_1_57_0 & i_2_1_135_0))))))) | (i_2_1_68_0 & ((~i_2_1_46_0 & i_2_1_135_0 & i_2_1_136_0) | (i_2_1_34_0 & (~i_2_1_46_0 | (~i_2_1_57_0 & i_2_1_135_0))))))) | ((i_2_1_135_0 | i_2_1_136_0) & ((i_2_1_34_0 & i_2_1_41_0 & ~i_2_1_57_0 & (~i_2_1_51_0 | i_2_1_68_0)) | (~i_2_1_46_0 & ~i_2_1_51_0 & i_2_1_68_0))) | (i_2_1_68_0 & ((i_2_1_136_0 & ((i_2_1_34_0 & i_2_1_135_0 & (i_2_1_41_0 | ~i_2_1_57_0)) | (i_2_1_41_0 & ~i_2_1_51_0 & ~i_2_1_57_0))) | (~i_2_1_57_0 & ((i_2_1_34_0 & (~i_2_1_46_0 | (~i_2_1_51_0 & i_2_1_135_0))) | (~i_2_1_46_0 & ~i_2_1_51_0))))) | (~i_2_1_46_0 & ~i_2_1_51_0 & (i_2_1_34_0 | (~i_2_1_57_0 & i_2_1_135_0 & i_2_1_136_0))))) | (i_2_1_41_0 & ((~i_2_1_51_0 & ((i_2_1_34_0 & i_2_1_68_0 & i_2_1_136_0) | (i_2_1_135_0 & ~i_2_1_136_0 & ~i_2_1_32_0 & ~i_2_1_46_0))) | (i_2_1_68_0 & ((i_2_1_135_0 & ((~i_2_1_46_0 & ~i_2_1_57_0) | (i_2_1_136_0 & ((~i_2_1_46_0 & i_2_1_70_0) | (i_2_1_34_0 & (~i_2_1_57_0 | i_2_1_70_0)))))) | (i_2_1_34_0 & ~i_2_1_46_0 & ~i_2_1_135_0))))) | (i_2_1_34_0 & ((i_2_1_68_0 & ((~i_2_1_51_0 & (~i_2_1_46_0 | (~i_2_1_57_0 & i_2_1_136_0))) | (~i_2_1_46_0 & i_2_1_70_0 & (~i_2_1_57_0 | i_2_1_135_0)))) | (i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_51_0 & i_2_1_70_0))) | (~i_2_1_57_0 & i_2_1_68_0 & i_2_1_70_0 & i_2_1_136_0 & (~i_2_1_46_0 | ~i_2_1_51_0)))) | (~i_2_1_57_0 & ((i_2_1_68_0 & ((~i_2_1_51_0 & ((~i_2_1_32_0 & ((i_2_1_70_0 & i_2_1_135_0 & ~i_2_1_136_0) | (i_2_1_41_0 & ~i_2_1_46_0))) | (i_2_1_34_0 & ((~i_2_1_49_0 & i_2_1_136_0) | (i_2_1_32_0 & i_2_1_41_0))) | (~i_2_1_49_0 & ((i_2_1_32_0 & ((~i_2_1_46_0 & i_2_1_70_0) | (i_2_1_41_0 & i_2_1_135_0 & i_2_1_136_0))) | (i_2_1_136_0 & ((~i_2_1_46_0 & i_2_1_135_0) | (i_2_1_41_0 & i_2_1_70_0))))) | (i_2_1_70_0 & i_2_1_135_0 & i_2_1_32_0 & i_2_1_41_0))) | (i_2_1_41_0 & ((i_2_1_136_0 & ((i_2_1_32_0 & i_2_1_34_0 & (~i_2_1_49_0 | ~i_2_1_135_0)) | (~i_2_1_46_0 & (i_2_1_70_0 | (~i_2_1_49_0 & ~i_2_1_135_0))))) | (~i_2_1_46_0 & ((~i_2_1_49_0 & i_2_1_70_0) | (i_2_1_32_0 & i_2_1_135_0))))) | (~i_2_1_46_0 & i_2_1_70_0 & ((~i_2_1_49_0 & (i_2_1_34_0 | i_2_1_135_0)) | (i_2_1_135_0 & (i_2_1_32_0 | i_2_1_136_0)))))) | (i_2_1_70_0 & ((i_2_1_136_0 & ((i_2_1_34_0 & (~i_2_1_41_0 | ~i_2_1_49_0)) | (~i_2_1_46_0 & ((i_2_1_41_0 & (~i_2_1_51_0 | (~i_2_1_49_0 & i_2_1_135_0))) | (i_2_1_32_0 & ~i_2_1_49_0 & ~i_2_1_51_0))) | (~i_2_1_38_0 & ~i_2_1_41_0 & ~i_2_1_49_0 & ~i_2_1_51_0 & i_2_1_135_0))) | (i_2_1_135_0 & ((i_2_1_32_0 & ((i_2_1_34_0 & (~i_2_1_46_0 | (~i_2_1_38_0 & ~i_2_1_51_0))) | (i_2_1_41_0 & (~i_2_1_46_0 | (~i_2_1_38_0 & ~i_2_1_49_0))))) | (i_2_1_34_0 & ~i_2_1_38_0 & ~i_2_1_49_0 & ~i_2_1_68_0))) | (i_2_1_34_0 & ~i_2_1_51_0 & ((~i_2_1_38_0 & ~i_2_1_46_0) | (i_2_1_32_0 & i_2_1_41_0 & ~i_2_1_136_0))))) | (~i_2_1_46_0 & ((i_2_1_34_0 & (i_2_1_136_0 | (~i_2_1_51_0 & i_2_1_135_0))) | (i_2_1_41_0 & ~i_2_1_49_0 & ~i_2_1_136_0 & (i_2_1_32_0 | (~i_2_1_70_0 & i_2_1_135_0))))))) | (~i_2_1_46_0 & ((i_2_1_41_0 & ((i_2_1_34_0 & ((i_2_1_68_0 & i_2_1_136_0) | (~i_2_1_49_0 & ~i_2_1_70_0))) | (i_2_1_32_0 & ((i_2_1_68_0 & ((~i_2_1_49_0 & (~i_2_1_51_0 | i_2_1_135_0)) | (~i_2_1_51_0 & i_2_1_70_0) | (i_2_1_51_0 & i_2_1_135_0 & i_2_1_136_0))) | (~i_2_1_49_0 & i_2_1_70_0 & i_2_1_135_0))) | (~i_2_1_49_0 & ~i_2_1_51_0 & i_2_1_136_0 & ((~i_2_1_70_0 & ~i_2_1_135_0) | (i_2_1_68_0 & i_2_1_70_0 & i_2_1_135_0))))) | (i_2_1_68_0 & ((i_2_1_34_0 & ((~i_2_1_49_0 & ~i_2_1_51_0 & i_2_1_135_0) | (i_2_1_32_0 & i_2_1_70_0 & ~i_2_1_135_0))) | (i_2_1_32_0 & ((~i_2_1_49_0 & ~i_2_1_51_0 & ((i_2_1_70_0 & i_2_1_135_0) | (i_2_1_57_0 & ~i_2_1_135_0 & i_2_1_136_0))) | (~i_2_1_135_0 & i_2_1_136_0 & i_2_1_47_0 & i_2_1_70_0))))) | (i_2_1_70_0 & i_2_1_136_0 & i_2_1_34_0 & ~i_2_1_51_0))) | (i_2_1_34_0 & ((~i_2_1_49_0 & ((i_2_1_68_0 & ((i_2_1_136_0 & ((i_2_1_41_0 & i_2_1_70_0 & i_2_1_135_0) | (i_2_1_32_0 & ~i_2_1_51_0 & (i_2_1_41_0 | ~i_2_1_135_0)))) | (i_2_1_32_0 & i_2_1_70_0 & i_2_1_135_0))) | (i_2_1_32_0 & ~i_2_1_38_0 & i_2_1_41_0 & ~i_2_1_51_0 & i_2_1_70_0))) | (i_2_1_70_0 & i_2_1_136_0 & i_2_1_32_0 & i_2_1_68_0))) | (i_2_1_32_0 & i_2_1_41_0 & ~i_2_1_49_0 & i_2_1_70_0 & i_2_1_136_0 & ~i_2_1_51_0 & i_2_1_68_0))) | (i_2_1_34_0 & ((i_2_1_32_0 & ((i_2_1_135_0 & ((i_2_1_70_0 & ((~i_2_1_13_0 & ((~i_2_1_57_0 & i_2_1_68_0) | (i_2_1_38_0 & ~i_2_1_51_0 & i_2_1_54_0 & i_2_1_57_0 & ~i_2_1_136_0))) | (~i_2_1_46_0 & ((i_2_1_38_0 & ~i_2_1_49_0) | (~i_2_1_38_0 & ~i_2_1_51_0 & ~i_2_1_57_0))) | (i_2_1_38_0 & ((~i_2_1_49_0 & ~i_2_1_51_0) | (i_2_1_41_0 & ~i_2_1_57_0 & i_2_1_136_0 & (~i_2_1_49_0 | ~i_2_1_51_0)))) | (i_2_1_41_0 & ~i_2_1_49_0 & ~i_2_1_51_0 & i_2_1_68_0 & i_2_1_136_0))) | (~i_2_1_46_0 & ((i_2_1_136_0 & ((~i_2_1_57_0 & i_2_1_68_0) | (~i_2_1_49_0 & i_2_1_51_0 & (i_2_1_47_0 | i_2_1_68_0)))) | (i_2_1_41_0 & i_2_1_68_0) | (~i_2_1_51_0 & ~i_2_1_57_0 & (i_2_1_68_0 | (i_2_1_38_0 & ~i_2_1_70_0))))) | (i_2_1_68_0 & ((i_2_1_38_0 & i_2_1_41_0 & ((~i_2_1_49_0 & i_2_1_136_0) | (i_2_1_49_0 & ~i_2_1_51_0 & ~i_2_1_136_0))) | (~i_2_1_57_0 & i_2_1_136_0 & ~i_2_1_49_0 & ~i_2_1_51_0))))) | (i_2_1_68_0 & ((i_2_1_38_0 & ((i_2_1_41_0 & ((i_2_1_57_0 & i_2_1_136_0 & (~i_2_1_49_0 | i_2_1_51_0)) | (~i_2_1_49_0 & ~i_2_1_57_0 & (~i_2_1_51_0 | i_2_1_70_0)))) | (~i_2_1_46_0 & ((~i_2_1_57_0 & ~i_2_1_136_0) | (~i_2_1_51_0 & (~i_2_1_49_0 | ~i_2_1_70_0)))) | (i_2_1_54_0 & i_2_1_70_0 & i_2_1_136_0))) | (~i_2_1_46_0 & ((~i_2_1_51_0 & ((i_2_1_41_0 & (~i_2_1_49_0 | i_2_1_70_0)) | (i_2_1_136_0 & (i_2_1_70_0 | (~i_2_1_49_0 & ~i_2_1_135_0))))) | (~i_2_1_57_0 & ((~i_2_1_49_0 & i_2_1_136_0) | (i_2_1_49_0 & i_2_1_70_0))))) | (~i_2_1_51_0 & ~i_2_1_57_0 & i_2_1_70_0))) | (~i_2_1_46_0 & ((~i_2_1_57_0 & ((~i_2_1_49_0 & ((i_2_1_41_0 & ~i_2_1_136_0) | (~i_2_1_41_0 & ~i_2_1_51_0))) | (i_2_1_41_0 & ((i_2_1_70_0 & i_2_1_136_0) | (~i_2_1_51_0 & ~i_2_1_136_0))))) | (i_2_1_38_0 & i_2_1_41_0 & ~i_2_1_49_0))))) | (~i_2_1_57_0 & ((~i_2_1_46_0 & ((~i_2_1_51_0 & ((~i_2_1_32_0 & ((i_2_1_38_0 & i_2_1_70_0 & i_2_1_135_0) | (~i_2_1_38_0 & ~i_2_1_70_0 & i_2_1_136_0))) | (i_2_1_68_0 & ((~i_2_1_49_0 & i_2_1_135_0) | (i_2_1_38_0 & i_2_1_49_0))))) | (i_2_1_68_0 & ((i_2_1_38_0 & ((i_2_1_135_0 & i_2_1_136_0) | (~i_2_1_49_0 & (i_2_1_136_0 | (i_2_1_41_0 & i_2_1_70_0))))) | (i_2_1_41_0 & (i_2_1_136_0 | (i_2_1_70_0 & i_2_1_135_0))) | (i_2_1_135_0 & i_2_1_136_0 & (~i_2_1_49_0 | i_2_1_70_0)))) | (i_2_1_41_0 & ~i_2_1_49_0 & i_2_1_135_0 & ((i_2_1_70_0 & i_2_1_136_0) | (~i_2_1_70_0 & ~i_2_1_136_0))))) | (i_2_1_68_0 & ((i_2_1_135_0 & ((i_2_1_38_0 & i_2_1_136_0 & ((~i_2_1_41_0 & i_2_1_70_0) | (i_2_1_41_0 & ~i_2_1_51_0))) | (~i_2_1_51_0 & i_2_1_70_0) | (i_2_1_41_0 & ~i_2_1_136_0 & ((~i_2_1_49_0 & i_2_1_70_0) | (i_2_1_49_0 & ~i_2_1_51_0))))) | (~i_2_1_49_0 & i_2_1_70_0 & (~i_2_1_51_0 | (i_2_1_38_0 & i_2_1_41_0 & i_2_1_136_0))))) | (i_2_1_38_0 & i_2_1_41_0 & ~i_2_1_49_0 & ~i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_51_0 & i_2_1_70_0))) | (i_2_1_68_0 & ((i_2_1_41_0 & ((~i_2_1_51_0 & ~i_2_1_135_0 & ((i_2_1_38_0 & i_2_1_70_0) | (~i_2_1_46_0 & i_2_1_136_0))) | (i_2_1_38_0 & ((~i_2_1_46_0 & ~i_2_1_49_0 & (i_2_1_135_0 | (i_2_1_70_0 & i_2_1_136_0))) | (i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0 & i_2_1_49_0 & i_2_1_57_0))) | (i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_46_0 & ~i_2_1_49_0))) | (i_2_1_38_0 & i_2_1_136_0 & ((~i_2_1_51_0 & i_2_1_70_0) | (~i_2_1_49_0 & i_2_1_135_0 & (~i_2_1_46_0 | (~i_2_1_41_0 & i_2_1_70_0))))))) | (i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0 & i_2_1_38_0 & ~i_2_1_46_0 & ~i_2_1_51_0))) | (i_2_1_68_0 & ((i_2_1_32_0 & ((i_2_1_38_0 & ((~i_2_1_51_0 & ((i_2_1_135_0 & ((~i_2_1_13_0 & i_2_1_49_0 & i_2_1_57_0 & (i_2_1_70_0 | (~i_2_1_41_0 & i_2_1_136_0))) | (i_2_1_70_0 & i_2_1_136_0) | (~i_2_1_57_0 & ((~i_2_1_49_0 & i_2_1_70_0) | (~i_2_1_41_0 & ~i_2_1_46_0))))) | (i_2_1_70_0 & ((i_2_1_41_0 & (~i_2_1_46_0 | (~i_2_1_49_0 & i_2_1_136_0))) | (~i_2_1_46_0 & ~i_2_1_57_0) | (i_2_1_49_0 & i_2_1_54_0 & i_2_1_57_0 & i_2_1_136_0))) | (~i_2_1_57_0 & i_2_1_136_0 & ~i_2_1_46_0 & i_2_1_49_0))) | (i_2_1_70_0 & ((~i_2_1_57_0 & ((i_2_1_41_0 & (~i_2_1_46_0 | (~i_2_1_49_0 & i_2_1_135_0 & i_2_1_136_0))) | (~i_2_1_46_0 & ~i_2_1_49_0 & i_2_1_136_0) | (i_2_1_135_0 & ~i_2_1_136_0 & ~i_2_1_41_0 & i_2_1_51_0))) | (i_2_1_135_0 & ((~i_2_1_41_0 & i_2_1_49_0 & i_2_1_57_0 & i_2_1_136_0) | (~i_2_1_46_0 & ~i_2_1_49_0 & i_2_1_51_0 & ~i_2_1_136_0))))) | (i_2_1_41_0 & ~i_2_1_46_0 & ((i_2_1_49_0 & i_2_1_57_0) | (~i_2_1_49_0 & i_2_1_135_0))))) | (i_2_1_41_0 & ~i_2_1_46_0 & ((~i_2_1_49_0 & ((~i_2_1_51_0 & ((~i_2_1_57_0 & i_2_1_136_0) | (i_2_1_70_0 & i_2_1_135_0))) | (i_2_1_51_0 & i_2_1_57_0 & i_2_1_70_0 & ~i_2_1_135_0 & i_2_1_136_0))) | (~i_2_1_57_0 & i_2_1_70_0 & (i_2_1_135_0 | (i_2_1_49_0 & i_2_1_136_0))))))) | (~i_2_1_46_0 & ((~i_2_1_49_0 & ((i_2_1_38_0 & ((i_2_1_41_0 & i_2_1_70_0 & (~i_2_1_51_0 | (~i_2_1_57_0 & i_2_1_135_0 & i_2_1_136_0))) | (~i_2_1_57_0 & i_2_1_135_0 & (~i_2_1_51_0 | (~i_2_1_32_0 & ~i_2_1_41_0 & ~i_2_1_70_0 & i_2_1_136_0))))) | (i_2_1_70_0 & i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_51_0 & ~i_2_1_57_0))) | (i_2_1_41_0 & ~i_2_1_51_0 & ~i_2_1_57_0 & i_2_1_70_0 & (i_2_1_135_0 | (i_2_1_49_0 & i_2_1_136_0))))) | (i_2_1_135_0 & i_2_1_136_0 & ~i_2_1_57_0 & i_2_1_70_0 & i_2_1_38_0 & ~i_2_1_49_0 & ~i_2_1_51_0))) | (i_2_1_32_0 & i_2_1_38_0 & ~i_2_1_46_0 & i_2_1_70_0 & ((i_2_1_41_0 & ((~i_2_1_51_0 & ~i_2_1_57_0 & i_2_1_135_0) | (~i_2_1_49_0 & i_2_1_136_0 & ((~i_2_1_57_0 & i_2_1_135_0) | (~i_2_1_51_0 & ~i_2_1_135_0))))) | (~i_2_1_49_0 & ~i_2_1_51_0 & ~i_2_1_57_0 & i_2_1_135_0 & ~i_2_1_136_0)));
endmodule
