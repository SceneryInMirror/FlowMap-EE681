// Benchmark "kernel_2_5" written by ABC on Wed May  4 16:43:15 2022

module kernel_2_5 ( 
    i_2_5_12_0, i_2_5_42_0, i_2_5_62_0, i_2_5_65_0, i_2_5_70_0, i_2_5_82_0,
    i_2_5_84_0, i_2_5_90_0, i_2_5_91_0, i_2_5_92_0, i_2_5_93_0, i_2_5_98_0,
    i_2_5_99_0, i_2_5_102_0, i_2_5_148_0,
    o_2_5_0_0  );
  input  i_2_5_12_0, i_2_5_42_0, i_2_5_62_0, i_2_5_65_0, i_2_5_70_0,
    i_2_5_82_0, i_2_5_84_0, i_2_5_90_0, i_2_5_91_0, i_2_5_92_0, i_2_5_93_0,
    i_2_5_98_0, i_2_5_99_0, i_2_5_102_0, i_2_5_148_0;
  output o_2_5_0_0;
  wire new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_,
    new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_,
    new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_,
    new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_;
  NOT      g0000(.a(i_2_5_92_0), .O(new_n17_));
  NOT      g0001(.a(i_2_5_93_0), .O(new_n18_));
  NOT      g0002(.a(i_2_5_98_0), .O(new_n19_));
  NOT      g0003(.a(i_2_5_99_0), .O(new_n20_));
  NOT      g0004(.a(i_2_5_90_0), .O(new_n21_));
  AND      g0005(.a(new_n21_), .b(i_2_5_84_0), .O(new_n22_));
  OR       g0006(.a(new_n22_), .b(i_2_5_82_0), .O(new_n23_));
  OR       g0007(.a(new_n21_), .b(i_2_5_84_0), .O(new_n24_));
  AND      g0008(.a(new_n24_), .b(i_2_5_12_0), .O(new_n25_));
  AND      g0009(.a(new_n25_), .b(new_n23_), .O(new_n26_));
  NOT      g0010(.a(i_2_5_65_0), .O(new_n27_));
  AND      g0011(.a(i_2_5_82_0), .b(i_2_5_12_0), .O(new_n28_));
  OR       g0012(.a(new_n28_), .b(new_n21_), .O(new_n29_));
  AND      g0013(.a(new_n29_), .b(new_n27_), .O(new_n30_));
  OR       g0014(.a(i_2_5_84_0), .b(i_2_5_12_0), .O(new_n31_));
  AND      g0015(.a(new_n31_), .b(new_n27_), .O(new_n32_));
  AND      g0016(.a(new_n21_), .b(i_2_5_82_0), .O(new_n33_));
  OR       g0017(.a(i_2_5_84_0), .b(new_n27_), .O(new_n34_));
  AND      g0018(.a(new_n34_), .b(new_n33_), .O(new_n35_));
  OR       g0019(.a(new_n35_), .b(new_n32_), .O(new_n36_));
  OR       g0020(.a(new_n36_), .b(new_n30_), .O(new_n37_));
  OR       g0021(.a(new_n37_), .b(new_n26_), .O(new_n38_));
  AND      g0022(.a(new_n38_), .b(i_2_5_62_0), .O(new_n39_));
  OR       g0023(.a(i_2_5_90_0), .b(i_2_5_65_0), .O(new_n40_));
  NOT      g0024(.a(new_n40_), .O(new_n41_));
  AND      g0025(.a(new_n41_), .b(new_n31_), .O(new_n42_));
  OR       g0026(.a(new_n42_), .b(new_n39_), .O(new_n43_));
  AND      g0027(.a(new_n43_), .b(i_2_5_102_0), .O(new_n44_));
  AND      g0028(.a(new_n27_), .b(i_2_5_62_0), .O(new_n45_));
  OR       g0029(.a(new_n45_), .b(new_n28_), .O(new_n46_));
  AND      g0030(.a(new_n46_), .b(new_n22_), .O(new_n47_));
  OR       g0031(.a(new_n47_), .b(new_n44_), .O(new_n48_));
  AND      g0032(.a(new_n48_), .b(new_n20_), .O(new_n49_));
  AND      g0033(.a(new_n27_), .b(i_2_5_12_0), .O(new_n50_));
  AND      g0034(.a(i_2_5_84_0), .b(new_n27_), .O(new_n51_));
  AND      g0035(.a(new_n51_), .b(i_2_5_102_0), .O(new_n52_));
  OR       g0036(.a(new_n52_), .b(new_n50_), .O(new_n53_));
  NOT      g0037(.a(i_2_5_91_0), .O(new_n54_));
  AND      g0038(.a(i_2_5_102_0), .b(new_n54_), .O(new_n55_));
  NAND     g0039(.a(i_2_5_102_0), .b(i_2_5_82_0), .O(new_n56_));
  NAND     g0040(.a(new_n56_), .b(i_2_5_99_0), .O(new_n57_));
  AND      g0041(.a(new_n57_), .b(i_2_5_84_0), .O(new_n58_));
  OR       g0042(.a(new_n58_), .b(new_n55_), .O(new_n59_));
  OR       g0043(.a(new_n59_), .b(new_n53_), .O(new_n60_));
  AND      g0044(.a(new_n60_), .b(i_2_5_62_0), .O(new_n61_));
  NOT      g0045(.a(i_2_5_62_0), .O(new_n62_));
  AND      g0046(.a(new_n56_), .b(i_2_5_91_0), .O(new_n63_));
  OR       g0047(.a(new_n63_), .b(new_n62_), .O(new_n64_));
  NOT      g0048(.a(i_2_5_102_0), .O(new_n65_));
  OR       g0049(.a(new_n65_), .b(i_2_5_99_0), .O(new_n66_));
  NOT      g0050(.a(i_2_5_70_0), .O(new_n67_));
  OR       g0051(.a(new_n67_), .b(i_2_5_65_0), .O(new_n68_));
  AND      g0052(.a(new_n68_), .b(new_n66_), .O(new_n69_));
  NAND     g0053(.a(new_n69_), .b(new_n64_), .O(new_n70_));
  AND      g0054(.a(new_n70_), .b(i_2_5_12_0), .O(new_n71_));
  OR       g0055(.a(i_2_5_102_0), .b(i_2_5_84_0), .O(new_n72_));
  AND      g0056(.a(new_n72_), .b(new_n54_), .O(new_n73_));
  OR       g0057(.a(i_2_5_102_0), .b(new_n27_), .O(new_n74_));
  AND      g0058(.a(new_n74_), .b(i_2_5_84_0), .O(new_n75_));
  OR       g0059(.a(new_n75_), .b(new_n20_), .O(new_n76_));
  AND      g0060(.a(new_n76_), .b(new_n73_), .O(new_n77_));
  AND      g0061(.a(i_2_5_82_0), .b(new_n27_), .O(new_n78_));
  AND      g0062(.a(new_n78_), .b(i_2_5_84_0), .O(new_n79_));
  OR       g0063(.a(new_n79_), .b(new_n77_), .O(new_n80_));
  OR       g0064(.a(new_n80_), .b(new_n71_), .O(new_n81_));
  OR       g0065(.a(new_n81_), .b(new_n61_), .O(new_n82_));
  AND      g0066(.a(new_n82_), .b(new_n21_), .O(new_n83_));
  OR       g0067(.a(i_2_5_99_0), .b(i_2_5_91_0), .O(new_n84_));
  NOT      g0068(.a(new_n84_), .O(new_n85_));
  NAND     g0069(.a(i_2_5_99_0), .b(i_2_5_91_0), .O(new_n86_));
  AND      g0070(.a(new_n86_), .b(new_n27_), .O(new_n87_));
  OR       g0071(.a(new_n87_), .b(new_n85_), .O(new_n88_));
  AND      g0072(.a(new_n88_), .b(i_2_5_82_0), .O(new_n89_));
  OR       g0073(.a(new_n27_), .b(i_2_5_12_0), .O(new_n90_));
  AND      g0074(.a(new_n90_), .b(new_n20_), .O(new_n91_));
  AND      g0075(.a(new_n54_), .b(i_2_5_82_0), .O(new_n92_));
  AND      g0076(.a(new_n92_), .b(new_n31_), .O(new_n93_));
  OR       g0077(.a(new_n93_), .b(new_n91_), .O(new_n94_));
  AND      g0078(.a(new_n94_), .b(i_2_5_62_0), .O(new_n95_));
  OR       g0079(.a(new_n95_), .b(new_n89_), .O(new_n96_));
  AND      g0080(.a(new_n96_), .b(i_2_5_102_0), .O(new_n97_));
  AND      g0081(.a(new_n90_), .b(new_n54_), .O(new_n98_));
  NOT      g0082(.a(i_2_5_42_0), .O(new_n99_));
  AND      g0083(.a(i_2_5_82_0), .b(new_n99_), .O(new_n100_));
  AND      g0084(.a(new_n100_), .b(new_n27_), .O(new_n101_));
  OR       g0085(.a(new_n101_), .b(new_n98_), .O(new_n102_));
  AND      g0086(.a(new_n102_), .b(i_2_5_102_0), .O(new_n103_));
  AND      g0087(.a(i_2_5_102_0), .b(new_n20_), .O(new_n104_));
  OR       g0088(.a(new_n104_), .b(new_n54_), .O(new_n105_));
  NAND     g0089(.a(i_2_5_99_0), .b(i_2_5_65_0), .O(new_n106_));
  AND      g0090(.a(new_n106_), .b(i_2_5_62_0), .O(new_n107_));
  AND      g0091(.a(new_n107_), .b(new_n105_), .O(new_n108_));
  OR       g0092(.a(new_n108_), .b(new_n103_), .O(new_n109_));
  AND      g0093(.a(new_n109_), .b(new_n24_), .O(new_n110_));
  NOT      g0094(.a(new_n45_), .O(new_n111_));
  NOT      g0095(.a(i_2_5_84_0), .O(new_n112_));
  OR       g0096(.a(new_n112_), .b(i_2_5_65_0), .O(new_n113_));
  OR       g0097(.a(new_n113_), .b(i_2_5_99_0), .O(new_n114_));
  NAND     g0098(.a(new_n114_), .b(new_n111_), .O(new_n115_));
  OR       g0099(.a(new_n54_), .b(i_2_5_84_0), .O(new_n116_));
  AND      g0100(.a(new_n116_), .b(new_n20_), .O(new_n117_));
  OR       g0101(.a(i_2_5_82_0), .b(i_2_5_42_0), .O(new_n118_));
  NAND     g0102(.a(new_n118_), .b(new_n62_), .O(new_n119_));
  AND      g0103(.a(new_n119_), .b(new_n117_), .O(new_n120_));
  AND      g0104(.a(new_n120_), .b(new_n115_), .O(new_n121_));
  AND      g0105(.a(new_n54_), .b(i_2_5_62_0), .O(new_n122_));
  OR       g0106(.a(new_n122_), .b(new_n20_), .O(new_n123_));
  AND      g0107(.a(i_2_5_84_0), .b(i_2_5_82_0), .O(new_n124_));
  OR       g0108(.a(new_n21_), .b(i_2_5_12_0), .O(new_n125_));
  AND      g0109(.a(new_n125_), .b(new_n124_), .O(new_n126_));
  OR       g0110(.a(new_n126_), .b(new_n50_), .O(new_n127_));
  AND      g0111(.a(new_n127_), .b(new_n123_), .O(new_n128_));
  OR       g0112(.a(i_2_5_102_0), .b(i_2_5_82_0), .O(new_n129_));
  NOT      g0113(.a(i_2_5_12_0), .O(new_n130_));
  OR       g0114(.a(new_n113_), .b(new_n130_), .O(new_n131_));
  OR       g0115(.a(new_n84_), .b(new_n62_), .O(new_n132_));
  NAND     g0116(.a(new_n132_), .b(new_n131_), .O(new_n133_));
  AND      g0117(.a(new_n133_), .b(new_n129_), .O(new_n134_));
  OR       g0118(.a(new_n134_), .b(new_n128_), .O(new_n135_));
  OR       g0119(.a(new_n135_), .b(new_n121_), .O(new_n136_));
  OR       g0120(.a(new_n136_), .b(new_n110_), .O(new_n137_));
  OR       g0121(.a(new_n137_), .b(new_n97_), .O(new_n138_));
  OR       g0122(.a(new_n138_), .b(new_n83_), .O(new_n139_));
  NAND     g0123(.a(new_n139_), .b(i_2_5_148_0), .O(new_n140_));
  OR       g0124(.a(i_2_5_90_0), .b(new_n112_), .O(new_n141_));
  OR       g0125(.a(new_n141_), .b(new_n65_), .O(new_n142_));
  NAND     g0126(.a(i_2_5_62_0), .b(i_2_5_12_0), .O(new_n143_));
  OR       g0127(.a(new_n143_), .b(i_2_5_65_0), .O(new_n144_));
  OR       g0128(.a(new_n144_), .b(new_n142_), .O(new_n145_));
  NAND     g0129(.a(new_n145_), .b(new_n140_), .O(new_n146_));
  OR       g0130(.a(new_n146_), .b(new_n49_), .O(new_n147_));
  OR       g0131(.a(i_2_5_102_0), .b(i_2_5_62_0), .O(new_n148_));
  AND      g0132(.a(new_n21_), .b(i_2_5_12_0), .O(new_n149_));
  OR       g0133(.a(new_n149_), .b(new_n20_), .O(new_n150_));
  AND      g0134(.a(new_n150_), .b(i_2_5_102_0), .O(new_n151_));
  OR       g0135(.a(new_n151_), .b(new_n91_), .O(new_n152_));
  AND      g0136(.a(new_n152_), .b(i_2_5_84_0), .O(new_n153_));
  OR       g0137(.a(i_2_5_99_0), .b(i_2_5_90_0), .O(new_n154_));
  NAND     g0138(.a(new_n154_), .b(new_n40_), .O(new_n155_));
  OR       g0139(.a(new_n155_), .b(new_n91_), .O(new_n156_));
  AND      g0140(.a(new_n156_), .b(i_2_5_102_0), .O(new_n157_));
  OR       g0141(.a(new_n157_), .b(new_n153_), .O(new_n158_));
  AND      g0142(.a(new_n158_), .b(i_2_5_62_0), .O(new_n159_));
  AND      g0143(.a(new_n28_), .b(new_n20_), .O(new_n160_));
  OR       g0144(.a(i_2_5_82_0), .b(i_2_5_12_0), .O(new_n161_));
  OR       g0145(.a(new_n161_), .b(new_n34_), .O(new_n162_));
  NAND     g0146(.a(new_n162_), .b(new_n20_), .O(new_n163_));
  NAND     g0147(.a(new_n163_), .b(new_n131_), .O(new_n164_));
  AND      g0148(.a(new_n164_), .b(new_n21_), .O(new_n165_));
  OR       g0149(.a(new_n165_), .b(new_n160_), .O(new_n166_));
  OR       g0150(.a(new_n166_), .b(new_n159_), .O(new_n167_));
  AND      g0151(.a(new_n167_), .b(new_n148_), .O(new_n168_));
  AND      g0152(.a(new_n72_), .b(new_n20_), .O(new_n169_));
  NAND     g0153(.a(i_2_5_102_0), .b(i_2_5_84_0), .O(new_n170_));
  NOT      g0154(.a(new_n170_), .O(new_n171_));
  AND      g0155(.a(new_n171_), .b(new_n125_), .O(new_n172_));
  OR       g0156(.a(new_n172_), .b(new_n169_), .O(new_n173_));
  AND      g0157(.a(new_n173_), .b(i_2_5_62_0), .O(new_n174_));
  AND      g0158(.a(i_2_5_102_0), .b(i_2_5_62_0), .O(new_n175_));
  OR       g0159(.a(new_n175_), .b(i_2_5_84_0), .O(new_n176_));
  AND      g0160(.a(new_n176_), .b(new_n149_), .O(new_n177_));
  AND      g0161(.a(i_2_5_84_0), .b(i_2_5_62_0), .O(new_n178_));
  NAND     g0162(.a(new_n178_), .b(new_n21_), .O(new_n179_));
  OR       g0163(.a(i_2_5_99_0), .b(i_2_5_42_0), .O(new_n180_));
  NAND     g0164(.a(new_n180_), .b(new_n179_), .O(new_n181_));
  AND      g0165(.a(new_n181_), .b(new_n27_), .O(new_n182_));
  OR       g0166(.a(new_n182_), .b(new_n177_), .O(new_n183_));
  OR       g0167(.a(new_n183_), .b(new_n174_), .O(new_n184_));
  AND      g0168(.a(new_n184_), .b(i_2_5_82_0), .O(new_n185_));
  OR       g0169(.a(i_2_5_102_0), .b(new_n21_), .O(new_n186_));
  NAND     g0170(.a(i_2_5_148_0), .b(i_2_5_84_0), .O(new_n187_));
  NAND     g0171(.a(new_n187_), .b(i_2_5_99_0), .O(new_n188_));
  AND      g0172(.a(new_n188_), .b(i_2_5_62_0), .O(new_n189_));
  OR       g0173(.a(i_2_5_148_0), .b(new_n27_), .O(new_n190_));
  AND      g0174(.a(new_n190_), .b(new_n20_), .O(new_n191_));
  OR       g0175(.a(new_n191_), .b(new_n189_), .O(new_n192_));
  AND      g0176(.a(new_n192_), .b(new_n186_), .O(new_n193_));
  NAND     g0177(.a(new_n170_), .b(i_2_5_99_0), .O(new_n194_));
  AND      g0178(.a(new_n194_), .b(new_n115_), .O(new_n195_));
  NOT      g0179(.a(new_n154_), .O(new_n196_));
  AND      g0180(.a(new_n196_), .b(new_n72_), .O(new_n197_));
  OR       g0181(.a(new_n27_), .b(i_2_5_62_0), .O(new_n198_));
  NOT      g0182(.a(i_2_5_148_0), .O(new_n199_));
  OR       g0183(.a(new_n199_), .b(i_2_5_99_0), .O(new_n200_));
  NAND     g0184(.a(new_n200_), .b(new_n142_), .O(new_n201_));
  AND      g0185(.a(new_n201_), .b(new_n198_), .O(new_n202_));
  OR       g0186(.a(new_n202_), .b(new_n197_), .O(new_n203_));
  OR       g0187(.a(new_n203_), .b(new_n195_), .O(new_n204_));
  OR       g0188(.a(new_n204_), .b(new_n193_), .O(new_n205_));
  AND      g0189(.a(new_n205_), .b(i_2_5_42_0), .O(new_n206_));
  OR       g0190(.a(new_n206_), .b(new_n185_), .O(new_n207_));
  OR       g0191(.a(new_n207_), .b(new_n168_), .O(new_n208_));
  AND      g0192(.a(new_n208_), .b(new_n54_), .O(new_n209_));
  AND      g0193(.a(new_n20_), .b(i_2_5_82_0), .O(new_n210_));
  NOT      g0194(.a(new_n210_), .O(new_n211_));
  OR       g0195(.a(i_2_5_91_0), .b(i_2_5_90_0), .O(new_n212_));
  NAND     g0196(.a(new_n212_), .b(new_n211_), .O(new_n213_));
  AND      g0197(.a(new_n213_), .b(new_n27_), .O(new_n214_));
  OR       g0198(.a(new_n178_), .b(i_2_5_82_0), .O(new_n215_));
  AND      g0199(.a(i_2_5_148_0), .b(new_n54_), .O(new_n216_));
  OR       g0200(.a(new_n216_), .b(new_n189_), .O(new_n217_));
  AND      g0201(.a(new_n217_), .b(new_n215_), .O(new_n218_));
  OR       g0202(.a(new_n218_), .b(new_n214_), .O(new_n219_));
  AND      g0203(.a(new_n219_), .b(i_2_5_102_0), .O(new_n220_));
  NOT      g0204(.a(i_2_5_82_0), .O(new_n221_));
  OR       g0205(.a(new_n65_), .b(i_2_5_65_0), .O(new_n222_));
  OR       g0206(.a(new_n222_), .b(new_n199_), .O(new_n223_));
  OR       g0207(.a(i_2_5_148_0), .b(i_2_5_102_0), .O(new_n224_));
  OR       g0208(.a(new_n224_), .b(new_n179_), .O(new_n225_));
  NAND     g0209(.a(new_n225_), .b(new_n223_), .O(new_n226_));
  AND      g0210(.a(new_n226_), .b(new_n221_), .O(new_n227_));
  OR       g0211(.a(new_n20_), .b(i_2_5_82_0), .O(new_n228_));
  NAND     g0212(.a(new_n228_), .b(new_n21_), .O(new_n229_));
  NAND     g0213(.a(new_n229_), .b(new_n200_), .O(new_n230_));
  AND      g0214(.a(new_n230_), .b(new_n54_), .O(new_n231_));
  OR       g0215(.a(new_n21_), .b(i_2_5_62_0), .O(new_n232_));
  AND      g0216(.a(new_n232_), .b(new_n216_), .O(new_n233_));
  OR       g0217(.a(i_2_5_91_0), .b(i_2_5_65_0), .O(new_n234_));
  NOT      g0218(.a(new_n234_), .O(new_n235_));
  OR       g0219(.a(new_n235_), .b(new_n78_), .O(new_n236_));
  OR       g0220(.a(new_n236_), .b(new_n233_), .O(new_n237_));
  AND      g0221(.a(new_n237_), .b(i_2_5_84_0), .O(new_n238_));
  OR       g0222(.a(new_n238_), .b(new_n231_), .O(new_n239_));
  OR       g0223(.a(new_n239_), .b(new_n227_), .O(new_n240_));
  OR       g0224(.a(new_n240_), .b(new_n220_), .O(new_n241_));
  AND      g0225(.a(new_n241_), .b(i_2_5_12_0), .O(new_n242_));
  NOT      g0226(.a(new_n223_), .O(new_n243_));
  AND      g0227(.a(new_n24_), .b(i_2_5_62_0), .O(new_n244_));
  OR       g0228(.a(new_n244_), .b(new_n22_), .O(new_n245_));
  AND      g0229(.a(new_n245_), .b(new_n243_), .O(new_n246_));
  AND      g0230(.a(new_n105_), .b(new_n27_), .O(new_n247_));
  OR       g0231(.a(i_2_5_148_0), .b(new_n21_), .O(new_n248_));
  AND      g0232(.a(new_n122_), .b(new_n21_), .O(new_n249_));
  AND      g0233(.a(new_n20_), .b(i_2_5_62_0), .O(new_n250_));
  OR       g0234(.a(new_n250_), .b(new_n55_), .O(new_n251_));
  OR       g0235(.a(new_n251_), .b(new_n249_), .O(new_n252_));
  AND      g0236(.a(new_n252_), .b(new_n248_), .O(new_n253_));
  OR       g0237(.a(new_n253_), .b(new_n247_), .O(new_n254_));
  AND      g0238(.a(new_n254_), .b(i_2_5_84_0), .O(new_n255_));
  OR       g0239(.a(new_n216_), .b(new_n104_), .O(new_n256_));
  OR       g0240(.a(new_n245_), .b(new_n45_), .O(new_n257_));
  AND      g0241(.a(new_n257_), .b(new_n256_), .O(new_n258_));
  OR       g0242(.a(new_n249_), .b(new_n233_), .O(new_n259_));
  AND      g0243(.a(new_n259_), .b(i_2_5_102_0), .O(new_n260_));
  AND      g0244(.a(i_2_5_148_0), .b(i_2_5_62_0), .O(new_n261_));
  AND      g0245(.a(new_n261_), .b(i_2_5_102_0), .O(new_n262_));
  OR       g0246(.a(new_n262_), .b(new_n41_), .O(new_n263_));
  AND      g0247(.a(new_n263_), .b(new_n20_), .O(new_n264_));
  OR       g0248(.a(new_n264_), .b(new_n260_), .O(new_n265_));
  OR       g0249(.a(new_n265_), .b(new_n258_), .O(new_n266_));
  OR       g0250(.a(new_n266_), .b(new_n255_), .O(new_n267_));
  AND      g0251(.a(new_n267_), .b(i_2_5_82_0), .O(new_n268_));
  OR       g0252(.a(new_n268_), .b(new_n246_), .O(new_n269_));
  OR       g0253(.a(new_n269_), .b(new_n242_), .O(new_n270_));
  AND      g0254(.a(new_n270_), .b(i_2_5_42_0), .O(new_n271_));
  OR       g0255(.a(new_n271_), .b(new_n209_), .O(new_n272_));
  OR       g0256(.a(new_n272_), .b(new_n147_), .O(new_n273_));
  AND      g0257(.a(new_n273_), .b(new_n19_), .O(new_n274_));
  AND      g0258(.a(new_n210_), .b(i_2_5_148_0), .O(new_n275_));
  NOT      g0259(.a(new_n187_), .O(new_n276_));
  OR       g0260(.a(i_2_5_99_0), .b(i_2_5_65_0), .O(new_n277_));
  NOT      g0261(.a(new_n277_), .O(new_n278_));
  NAND     g0262(.a(i_2_5_84_0), .b(i_2_5_42_0), .O(new_n279_));
  NAND     g0263(.a(new_n279_), .b(i_2_5_99_0), .O(new_n280_));
  AND      g0264(.a(new_n280_), .b(i_2_5_82_0), .O(new_n281_));
  OR       g0265(.a(new_n281_), .b(new_n278_), .O(new_n282_));
  OR       g0266(.a(new_n282_), .b(new_n276_), .O(new_n283_));
  AND      g0267(.a(new_n283_), .b(new_n54_), .O(new_n284_));
  OR       g0268(.a(new_n284_), .b(new_n275_), .O(new_n285_));
  AND      g0269(.a(new_n285_), .b(new_n148_), .O(new_n286_));
  AND      g0270(.a(i_2_5_84_0), .b(new_n221_), .O(new_n287_));
  OR       g0271(.a(new_n287_), .b(new_n92_), .O(new_n288_));
  AND      g0272(.a(new_n288_), .b(i_2_5_42_0), .O(new_n289_));
  OR       g0273(.a(new_n289_), .b(new_n88_), .O(new_n290_));
  AND      g0274(.a(new_n290_), .b(i_2_5_102_0), .O(new_n291_));
  AND      g0275(.a(new_n92_), .b(new_n34_), .O(new_n292_));
  OR       g0276(.a(new_n292_), .b(new_n291_), .O(new_n293_));
  AND      g0277(.a(new_n293_), .b(i_2_5_148_0), .O(new_n294_));
  AND      g0278(.a(new_n54_), .b(i_2_5_84_0), .O(new_n295_));
  AND      g0279(.a(new_n295_), .b(new_n278_), .O(new_n296_));
  OR       g0280(.a(i_2_5_148_0), .b(new_n54_), .O(new_n297_));
  AND      g0281(.a(new_n27_), .b(i_2_5_42_0), .O(new_n298_));
  AND      g0282(.a(new_n298_), .b(new_n57_), .O(new_n299_));
  AND      g0283(.a(new_n124_), .b(i_2_5_102_0), .O(new_n300_));
  AND      g0284(.a(new_n300_), .b(i_2_5_62_0), .O(new_n301_));
  OR       g0285(.a(new_n301_), .b(new_n299_), .O(new_n302_));
  AND      g0286(.a(new_n302_), .b(new_n297_), .O(new_n303_));
  OR       g0287(.a(new_n303_), .b(new_n296_), .O(new_n304_));
  OR       g0288(.a(new_n304_), .b(new_n294_), .O(new_n305_));
  OR       g0289(.a(new_n78_), .b(i_2_5_42_0), .O(new_n306_));
  AND      g0290(.a(new_n306_), .b(i_2_5_62_0), .O(new_n307_));
  OR       g0291(.a(new_n250_), .b(new_n85_), .O(new_n308_));
  OR       g0292(.a(new_n308_), .b(new_n235_), .O(new_n309_));
  OR       g0293(.a(new_n309_), .b(new_n307_), .O(new_n310_));
  AND      g0294(.a(new_n310_), .b(new_n31_), .O(new_n311_));
  AND      g0295(.a(new_n88_), .b(i_2_5_62_0), .O(new_n312_));
  AND      g0296(.a(new_n54_), .b(i_2_5_42_0), .O(new_n313_));
  OR       g0297(.a(new_n313_), .b(new_n78_), .O(new_n314_));
  AND      g0298(.a(new_n314_), .b(new_n20_), .O(new_n315_));
  OR       g0299(.a(new_n315_), .b(new_n312_), .O(new_n316_));
  OR       g0300(.a(new_n316_), .b(new_n311_), .O(new_n317_));
  AND      g0301(.a(new_n317_), .b(new_n224_), .O(new_n318_));
  AND      g0302(.a(i_2_5_82_0), .b(i_2_5_42_0), .O(new_n319_));
  AND      g0303(.a(new_n319_), .b(i_2_5_102_0), .O(new_n320_));
  OR       g0304(.a(new_n320_), .b(new_n51_), .O(new_n321_));
  AND      g0305(.a(new_n321_), .b(new_n86_), .O(new_n322_));
  OR       g0306(.a(i_2_5_84_0), .b(i_2_5_42_0), .O(new_n323_));
  NAND     g0307(.a(new_n223_), .b(new_n84_), .O(new_n324_));
  AND      g0308(.a(new_n324_), .b(new_n323_), .O(new_n325_));
  OR       g0309(.a(new_n221_), .b(i_2_5_65_0), .O(new_n326_));
  NAND     g0310(.a(i_2_5_148_0), .b(i_2_5_102_0), .O(new_n327_));
  AND      g0311(.a(new_n327_), .b(i_2_5_99_0), .O(new_n328_));
  OR       g0312(.a(new_n328_), .b(new_n326_), .O(new_n329_));
  NAND     g0313(.a(new_n55_), .b(i_2_5_148_0), .O(new_n330_));
  NAND     g0314(.a(new_n330_), .b(new_n329_), .O(new_n331_));
  OR       g0315(.a(new_n331_), .b(new_n325_), .O(new_n332_));
  OR       g0316(.a(new_n332_), .b(new_n322_), .O(new_n333_));
  AND      g0317(.a(new_n333_), .b(i_2_5_62_0), .O(new_n334_));
  OR       g0318(.a(new_n334_), .b(new_n318_), .O(new_n335_));
  OR       g0319(.a(new_n335_), .b(new_n305_), .O(new_n336_));
  OR       g0320(.a(new_n336_), .b(new_n286_), .O(new_n337_));
  NAND     g0321(.a(i_2_5_148_0), .b(i_2_5_82_0), .O(new_n338_));
  NAND     g0322(.a(new_n338_), .b(i_2_5_99_0), .O(new_n339_));
  AND      g0323(.a(new_n339_), .b(i_2_5_102_0), .O(new_n340_));
  AND      g0324(.a(new_n261_), .b(i_2_5_84_0), .O(new_n341_));
  OR       g0325(.a(new_n341_), .b(new_n340_), .O(new_n342_));
  NAND     g0326(.a(new_n327_), .b(i_2_5_91_0), .O(new_n343_));
  AND      g0327(.a(new_n343_), .b(i_2_5_62_0), .O(new_n344_));
  NAND     g0328(.a(new_n170_), .b(i_2_5_91_0), .O(new_n345_));
  AND      g0329(.a(new_n345_), .b(new_n194_), .O(new_n346_));
  OR       g0330(.a(new_n346_), .b(new_n344_), .O(new_n347_));
  OR       g0331(.a(new_n347_), .b(new_n342_), .O(new_n348_));
  AND      g0332(.a(new_n348_), .b(new_n27_), .O(new_n349_));
  AND      g0333(.a(new_n116_), .b(i_2_5_148_0), .O(new_n350_));
  NOT      g0334(.a(new_n338_), .O(new_n351_));
  OR       g0335(.a(i_2_5_84_0), .b(i_2_5_82_0), .O(new_n352_));
  AND      g0336(.a(new_n352_), .b(new_n54_), .O(new_n353_));
  OR       g0337(.a(new_n353_), .b(new_n351_), .O(new_n354_));
  AND      g0338(.a(new_n354_), .b(i_2_5_62_0), .O(new_n355_));
  OR       g0339(.a(new_n355_), .b(new_n350_), .O(new_n356_));
  AND      g0340(.a(new_n356_), .b(i_2_5_102_0), .O(new_n357_));
  OR       g0341(.a(new_n326_), .b(i_2_5_148_0), .O(new_n358_));
  OR       g0342(.a(new_n358_), .b(new_n148_), .O(new_n359_));
  AND      g0343(.a(new_n187_), .b(new_n84_), .O(new_n360_));
  NAND     g0344(.a(new_n360_), .b(new_n359_), .O(new_n361_));
  AND      g0345(.a(new_n361_), .b(i_2_5_42_0), .O(new_n362_));
  NAND     g0346(.a(i_2_5_91_0), .b(i_2_5_65_0), .O(new_n363_));
  OR       g0347(.a(new_n250_), .b(new_n124_), .O(new_n364_));
  AND      g0348(.a(new_n364_), .b(new_n363_), .O(new_n365_));
  AND      g0349(.a(new_n122_), .b(i_2_5_148_0), .O(new_n366_));
  OR       g0350(.a(i_2_5_148_0), .b(new_n20_), .O(new_n367_));
  AND      g0351(.a(new_n367_), .b(new_n124_), .O(new_n368_));
  OR       g0352(.a(new_n368_), .b(new_n366_), .O(new_n369_));
  OR       g0353(.a(new_n369_), .b(new_n365_), .O(new_n370_));
  OR       g0354(.a(new_n370_), .b(new_n362_), .O(new_n371_));
  OR       g0355(.a(new_n371_), .b(new_n357_), .O(new_n372_));
  OR       g0356(.a(new_n372_), .b(new_n349_), .O(new_n373_));
  AND      g0357(.a(new_n373_), .b(i_2_5_12_0), .O(new_n374_));
  OR       g0358(.a(new_n313_), .b(new_n27_), .O(new_n375_));
  AND      g0359(.a(new_n375_), .b(i_2_5_84_0), .O(new_n376_));
  OR       g0360(.a(new_n178_), .b(i_2_5_12_0), .O(new_n377_));
  OR       g0361(.a(new_n175_), .b(i_2_5_148_0), .O(new_n378_));
  AND      g0362(.a(new_n378_), .b(new_n377_), .O(new_n379_));
  AND      g0363(.a(i_2_5_62_0), .b(i_2_5_42_0), .O(new_n380_));
  OR       g0364(.a(i_2_5_148_0), .b(i_2_5_84_0), .O(new_n381_));
  NOT      g0365(.a(new_n381_), .O(new_n382_));
  AND      g0366(.a(new_n382_), .b(new_n380_), .O(new_n383_));
  OR       g0367(.a(new_n383_), .b(new_n216_), .O(new_n384_));
  OR       g0368(.a(new_n384_), .b(new_n379_), .O(new_n385_));
  OR       g0369(.a(new_n385_), .b(new_n376_), .O(new_n386_));
  AND      g0370(.a(new_n386_), .b(i_2_5_82_0), .O(new_n387_));
  OR       g0371(.a(new_n178_), .b(new_n54_), .O(new_n388_));
  OR       g0372(.a(i_2_5_102_0), .b(i_2_5_12_0), .O(new_n389_));
  OR       g0373(.a(new_n389_), .b(i_2_5_148_0), .O(new_n390_));
  AND      g0374(.a(new_n390_), .b(new_n388_), .O(new_n391_));
  OR       g0375(.a(i_2_5_84_0), .b(i_2_5_62_0), .O(new_n392_));
  AND      g0376(.a(new_n392_), .b(new_n54_), .O(new_n393_));
  OR       g0377(.a(new_n393_), .b(new_n308_), .O(new_n394_));
  OR       g0378(.a(new_n394_), .b(new_n391_), .O(new_n395_));
  AND      g0379(.a(new_n395_), .b(new_n27_), .O(new_n396_));
  AND      g0380(.a(new_n20_), .b(i_2_5_12_0), .O(new_n397_));
  OR       g0381(.a(new_n397_), .b(new_n148_), .O(new_n398_));
  AND      g0382(.a(new_n367_), .b(new_n54_), .O(new_n399_));
  AND      g0383(.a(new_n399_), .b(new_n398_), .O(new_n400_));
  OR       g0384(.a(new_n250_), .b(new_n276_), .O(new_n401_));
  AND      g0385(.a(new_n401_), .b(i_2_5_102_0), .O(new_n402_));
  OR       g0386(.a(new_n85_), .b(new_n51_), .O(new_n403_));
  AND      g0387(.a(new_n403_), .b(i_2_5_42_0), .O(new_n404_));
  OR       g0388(.a(new_n404_), .b(new_n402_), .O(new_n405_));
  OR       g0389(.a(new_n405_), .b(new_n400_), .O(new_n406_));
  OR       g0390(.a(i_2_5_99_0), .b(new_n112_), .O(new_n407_));
  OR       g0391(.a(new_n198_), .b(new_n56_), .O(new_n408_));
  NAND     g0392(.a(new_n408_), .b(new_n407_), .O(new_n409_));
  AND      g0393(.a(new_n409_), .b(new_n99_), .O(new_n410_));
  AND      g0394(.a(new_n224_), .b(new_n54_), .O(new_n411_));
  OR       g0395(.a(new_n411_), .b(i_2_5_62_0), .O(new_n412_));
  AND      g0396(.a(new_n86_), .b(new_n31_), .O(new_n413_));
  AND      g0397(.a(new_n413_), .b(new_n412_), .O(new_n414_));
  OR       g0398(.a(new_n414_), .b(new_n410_), .O(new_n415_));
  OR       g0399(.a(new_n415_), .b(new_n406_), .O(new_n416_));
  OR       g0400(.a(new_n416_), .b(new_n396_), .O(new_n417_));
  OR       g0401(.a(new_n417_), .b(new_n387_), .O(new_n418_));
  AND      g0402(.a(new_n418_), .b(new_n21_), .O(new_n419_));
  OR       g0403(.a(new_n419_), .b(new_n374_), .O(new_n420_));
  OR       g0404(.a(new_n420_), .b(new_n337_), .O(new_n421_));
  AND      g0405(.a(new_n421_), .b(new_n19_), .O(new_n422_));
  AND      g0406(.a(new_n72_), .b(i_2_5_82_0), .O(new_n423_));
  OR       g0407(.a(new_n423_), .b(new_n345_), .O(new_n424_));
  AND      g0408(.a(new_n424_), .b(new_n27_), .O(new_n425_));
  AND      g0409(.a(i_2_5_102_0), .b(i_2_5_42_0), .O(new_n426_));
  OR       g0410(.a(new_n426_), .b(new_n117_), .O(new_n427_));
  OR       g0411(.a(new_n427_), .b(new_n425_), .O(new_n428_));
  AND      g0412(.a(new_n428_), .b(i_2_5_12_0), .O(new_n429_));
  OR       g0413(.a(new_n298_), .b(new_n55_), .O(new_n430_));
  AND      g0414(.a(new_n430_), .b(new_n20_), .O(new_n431_));
  NOT      g0415(.a(new_n279_), .O(new_n432_));
  AND      g0416(.a(new_n432_), .b(i_2_5_102_0), .O(new_n433_));
  OR       g0417(.a(new_n433_), .b(i_2_5_82_0), .O(new_n434_));
  AND      g0418(.a(new_n323_), .b(i_2_5_102_0), .O(new_n435_));
  AND      g0419(.a(new_n435_), .b(new_n375_), .O(new_n436_));
  AND      g0420(.a(new_n295_), .b(i_2_5_42_0), .O(new_n437_));
  OR       g0421(.a(new_n437_), .b(new_n221_), .O(new_n438_));
  OR       g0422(.a(new_n438_), .b(new_n436_), .O(new_n439_));
  AND      g0423(.a(new_n439_), .b(new_n434_), .O(new_n440_));
  OR       g0424(.a(new_n440_), .b(new_n431_), .O(new_n441_));
  OR       g0425(.a(new_n441_), .b(new_n429_), .O(new_n442_));
  AND      g0426(.a(new_n442_), .b(i_2_5_148_0), .O(new_n443_));
  AND      g0427(.a(i_2_5_84_0), .b(i_2_5_12_0), .O(new_n444_));
  AND      g0428(.a(new_n34_), .b(i_2_5_42_0), .O(new_n445_));
  OR       g0429(.a(new_n445_), .b(new_n444_), .O(new_n446_));
  AND      g0430(.a(new_n446_), .b(i_2_5_82_0), .O(new_n447_));
  AND      g0431(.a(new_n90_), .b(i_2_5_102_0), .O(new_n448_));
  AND      g0432(.a(new_n448_), .b(new_n447_), .O(new_n449_));
  AND      g0433(.a(new_n72_), .b(new_n27_), .O(new_n450_));
  OR       g0434(.a(new_n450_), .b(new_n118_), .O(new_n451_));
  AND      g0435(.a(new_n74_), .b(new_n20_), .O(new_n452_));
  AND      g0436(.a(new_n452_), .b(new_n451_), .O(new_n453_));
  OR       g0437(.a(new_n453_), .b(new_n449_), .O(new_n454_));
  AND      g0438(.a(new_n454_), .b(new_n54_), .O(new_n455_));
  NAND     g0439(.a(new_n161_), .b(new_n20_), .O(new_n456_));
  NOT      g0440(.a(new_n456_), .O(new_n457_));
  AND      g0441(.a(i_2_5_42_0), .b(i_2_5_12_0), .O(new_n458_));
  NAND     g0442(.a(new_n458_), .b(i_2_5_82_0), .O(new_n459_));
  NAND     g0443(.a(new_n459_), .b(new_n222_), .O(new_n460_));
  AND      g0444(.a(new_n460_), .b(new_n457_), .O(new_n461_));
  OR       g0445(.a(new_n461_), .b(new_n455_), .O(new_n462_));
  OR       g0446(.a(new_n462_), .b(new_n443_), .O(new_n463_));
  AND      g0447(.a(new_n463_), .b(i_2_5_62_0), .O(new_n464_));
  AND      g0448(.a(new_n458_), .b(i_2_5_84_0), .O(new_n465_));
  AND      g0449(.a(new_n31_), .b(i_2_5_102_0), .O(new_n466_));
  AND      g0450(.a(new_n466_), .b(new_n54_), .O(new_n467_));
  OR       g0451(.a(new_n467_), .b(new_n465_), .O(new_n468_));
  NAND     g0452(.a(new_n468_), .b(i_2_5_62_0), .O(new_n469_));
  AND      g0453(.a(i_2_5_102_0), .b(i_2_5_12_0), .O(new_n470_));
  NAND     g0454(.a(new_n470_), .b(new_n124_), .O(new_n471_));
  NAND     g0455(.a(new_n471_), .b(new_n469_), .O(new_n472_));
  AND      g0456(.a(new_n472_), .b(new_n367_), .O(new_n473_));
  NOT      g0457(.a(new_n319_), .O(new_n474_));
  AND      g0458(.a(new_n352_), .b(new_n228_), .O(new_n475_));
  NAND     g0459(.a(new_n475_), .b(new_n188_), .O(new_n476_));
  NAND     g0460(.a(new_n476_), .b(new_n474_), .O(new_n477_));
  AND      g0461(.a(new_n477_), .b(new_n54_), .O(new_n478_));
  NAND     g0462(.a(new_n407_), .b(new_n330_), .O(new_n479_));
  AND      g0463(.a(new_n479_), .b(new_n27_), .O(new_n480_));
  OR       g0464(.a(new_n319_), .b(i_2_5_148_0), .O(new_n481_));
  OR       g0465(.a(new_n481_), .b(new_n313_), .O(new_n482_));
  AND      g0466(.a(new_n482_), .b(new_n104_), .O(new_n483_));
  OR       g0467(.a(new_n483_), .b(new_n480_), .O(new_n484_));
  OR       g0468(.a(new_n484_), .b(new_n478_), .O(new_n485_));
  AND      g0469(.a(new_n485_), .b(i_2_5_12_0), .O(new_n486_));
  AND      g0470(.a(new_n326_), .b(new_n65_), .O(new_n487_));
  OR       g0471(.a(i_2_5_91_0), .b(new_n99_), .O(new_n488_));
  AND      g0472(.a(new_n488_), .b(i_2_5_99_0), .O(new_n489_));
  OR       g0473(.a(new_n489_), .b(new_n199_), .O(new_n490_));
  OR       g0474(.a(new_n490_), .b(new_n487_), .O(new_n491_));
  OR       g0475(.a(new_n92_), .b(i_2_5_42_0), .O(new_n492_));
  NAND     g0476(.a(new_n56_), .b(i_2_5_91_0), .O(new_n493_));
  AND      g0477(.a(new_n493_), .b(new_n20_), .O(new_n494_));
  NAND     g0478(.a(new_n494_), .b(new_n492_), .O(new_n495_));
  NAND     g0479(.a(new_n495_), .b(new_n491_), .O(new_n496_));
  AND      g0480(.a(new_n496_), .b(i_2_5_84_0), .O(new_n497_));
  AND      g0481(.a(i_2_5_102_0), .b(i_2_5_90_0), .O(new_n498_));
  AND      g0482(.a(i_2_5_148_0), .b(new_n20_), .O(new_n499_));
  OR       g0483(.a(new_n21_), .b(i_2_5_42_0), .O(new_n500_));
  AND      g0484(.a(new_n500_), .b(new_n499_), .O(new_n501_));
  AND      g0485(.a(new_n501_), .b(new_n498_), .O(new_n502_));
  AND      g0486(.a(new_n57_), .b(i_2_5_148_0), .O(new_n503_));
  AND      g0487(.a(new_n129_), .b(i_2_5_42_0), .O(new_n504_));
  AND      g0488(.a(new_n504_), .b(new_n20_), .O(new_n505_));
  OR       g0489(.a(new_n505_), .b(new_n503_), .O(new_n506_));
  AND      g0490(.a(new_n506_), .b(new_n235_), .O(new_n507_));
  OR       g0491(.a(new_n507_), .b(new_n502_), .O(new_n508_));
  OR       g0492(.a(new_n508_), .b(new_n497_), .O(new_n509_));
  OR       g0493(.a(new_n509_), .b(new_n486_), .O(new_n510_));
  OR       g0494(.a(new_n510_), .b(new_n473_), .O(new_n511_));
  OR       g0495(.a(new_n511_), .b(new_n464_), .O(new_n512_));
  OR       g0496(.a(new_n512_), .b(new_n422_), .O(new_n513_));
  AND      g0497(.a(new_n513_), .b(new_n67_), .O(new_n514_));
  OR       g0498(.a(new_n381_), .b(new_n67_), .O(new_n515_));
  AND      g0499(.a(new_n515_), .b(new_n104_), .O(new_n516_));
  AND      g0500(.a(new_n194_), .b(new_n67_), .O(new_n517_));
  OR       g0501(.a(new_n112_), .b(i_2_5_70_0), .O(new_n518_));
  OR       g0502(.a(new_n518_), .b(new_n199_), .O(new_n519_));
  OR       g0503(.a(new_n170_), .b(new_n199_), .O(new_n520_));
  NAND     g0504(.a(new_n520_), .b(new_n519_), .O(new_n521_));
  OR       g0505(.a(new_n521_), .b(new_n517_), .O(new_n522_));
  AND      g0506(.a(new_n522_), .b(i_2_5_82_0), .O(new_n523_));
  OR       g0507(.a(new_n523_), .b(new_n516_), .O(new_n524_));
  AND      g0508(.a(new_n524_), .b(new_n54_), .O(new_n525_));
  OR       g0509(.a(new_n221_), .b(i_2_5_70_0), .O(new_n526_));
  NOT      g0510(.a(new_n526_), .O(new_n527_));
  AND      g0511(.a(new_n527_), .b(new_n104_), .O(new_n528_));
  OR       g0512(.a(i_2_5_91_0), .b(i_2_5_84_0), .O(new_n529_));
  OR       g0513(.a(new_n529_), .b(i_2_5_65_0), .O(new_n530_));
  NAND     g0514(.a(new_n530_), .b(new_n187_), .O(new_n531_));
  AND      g0515(.a(new_n531_), .b(i_2_5_82_0), .O(new_n532_));
  AND      g0516(.a(new_n297_), .b(new_n67_), .O(new_n533_));
  OR       g0517(.a(i_2_5_148_0), .b(i_2_5_82_0), .O(new_n534_));
  NOT      g0518(.a(new_n534_), .O(new_n535_));
  AND      g0519(.a(i_2_5_102_0), .b(new_n112_), .O(new_n536_));
  AND      g0520(.a(new_n536_), .b(new_n535_), .O(new_n537_));
  OR       g0521(.a(new_n537_), .b(new_n533_), .O(new_n538_));
  AND      g0522(.a(new_n538_), .b(i_2_5_62_0), .O(new_n539_));
  AND      g0523(.a(new_n424_), .b(new_n104_), .O(new_n540_));
  OR       g0524(.a(new_n540_), .b(new_n539_), .O(new_n541_));
  OR       g0525(.a(new_n541_), .b(new_n532_), .O(new_n542_));
  AND      g0526(.a(new_n542_), .b(i_2_5_12_0), .O(new_n543_));
  OR       g0527(.a(new_n543_), .b(new_n528_), .O(new_n544_));
  OR       g0528(.a(new_n544_), .b(new_n525_), .O(new_n545_));
  NAND     g0529(.a(i_2_5_99_0), .b(i_2_5_84_0), .O(new_n546_));
  AND      g0530(.a(new_n546_), .b(new_n73_), .O(new_n547_));
  OR       g0531(.a(new_n547_), .b(new_n216_), .O(new_n548_));
  AND      g0532(.a(new_n548_), .b(new_n194_), .O(new_n549_));
  OR       g0533(.a(i_2_5_102_0), .b(new_n112_), .O(new_n550_));
  OR       g0534(.a(i_2_5_148_0), .b(new_n221_), .O(new_n551_));
  OR       g0535(.a(new_n551_), .b(new_n550_), .O(new_n552_));
  OR       g0536(.a(new_n552_), .b(new_n19_), .O(new_n553_));
  NAND     g0537(.a(new_n553_), .b(new_n84_), .O(new_n554_));
  AND      g0538(.a(new_n554_), .b(new_n67_), .O(new_n555_));
  OR       g0539(.a(new_n73_), .b(new_n20_), .O(new_n556_));
  OR       g0540(.a(new_n351_), .b(new_n300_), .O(new_n557_));
  AND      g0541(.a(new_n557_), .b(new_n556_), .O(new_n558_));
  OR       g0542(.a(new_n558_), .b(new_n555_), .O(new_n559_));
  OR       g0543(.a(new_n559_), .b(new_n549_), .O(new_n560_));
  AND      g0544(.a(new_n560_), .b(i_2_5_62_0), .O(new_n561_));
  AND      g0545(.a(new_n199_), .b(i_2_5_84_0), .O(new_n562_));
  NOT      g0546(.a(new_n327_), .O(new_n563_));
  OR       g0547(.a(new_n563_), .b(new_n122_), .O(new_n564_));
  OR       g0548(.a(new_n564_), .b(new_n562_), .O(new_n565_));
  NAND     g0549(.a(new_n381_), .b(i_2_5_82_0), .O(new_n566_));
  NAND     g0550(.a(new_n566_), .b(new_n56_), .O(new_n567_));
  NAND     g0551(.a(i_2_5_102_0), .b(i_2_5_91_0), .O(new_n568_));
  AND      g0552(.a(new_n568_), .b(new_n148_), .O(new_n569_));
  OR       g0553(.a(new_n569_), .b(new_n67_), .O(new_n570_));
  AND      g0554(.a(new_n570_), .b(new_n567_), .O(new_n571_));
  AND      g0555(.a(new_n571_), .b(new_n565_), .O(new_n572_));
  OR       g0556(.a(new_n518_), .b(i_2_5_12_0), .O(new_n573_));
  NAND     g0557(.a(new_n573_), .b(new_n84_), .O(new_n574_));
  AND      g0558(.a(new_n574_), .b(i_2_5_62_0), .O(new_n575_));
  AND      g0559(.a(new_n346_), .b(new_n67_), .O(new_n576_));
  AND      g0560(.a(i_2_5_102_0), .b(new_n67_), .O(new_n577_));
  OR       g0561(.a(new_n577_), .b(new_n276_), .O(new_n578_));
  AND      g0562(.a(new_n221_), .b(i_2_5_62_0), .O(new_n579_));
  OR       g0563(.a(new_n579_), .b(new_n92_), .O(new_n580_));
  AND      g0564(.a(new_n580_), .b(new_n578_), .O(new_n581_));
  AND      g0565(.a(new_n85_), .b(i_2_5_102_0), .O(new_n582_));
  OR       g0566(.a(new_n582_), .b(new_n581_), .O(new_n583_));
  OR       g0567(.a(new_n583_), .b(new_n576_), .O(new_n584_));
  OR       g0568(.a(new_n584_), .b(new_n575_), .O(new_n585_));
  OR       g0569(.a(new_n585_), .b(new_n572_), .O(new_n586_));
  AND      g0570(.a(new_n586_), .b(new_n27_), .O(new_n587_));
  OR       g0571(.a(new_n587_), .b(new_n561_), .O(new_n588_));
  OR       g0572(.a(new_n588_), .b(new_n545_), .O(new_n589_));
  AND      g0573(.a(new_n589_), .b(i_2_5_42_0), .O(new_n590_));
  OR       g0574(.a(new_n235_), .b(new_n51_), .O(new_n591_));
  OR       g0575(.a(new_n591_), .b(new_n73_), .O(new_n592_));
  AND      g0576(.a(new_n592_), .b(i_2_5_62_0), .O(new_n593_));
  OR       g0577(.a(new_n55_), .b(new_n27_), .O(new_n594_));
  AND      g0578(.a(new_n594_), .b(i_2_5_82_0), .O(new_n595_));
  AND      g0579(.a(new_n222_), .b(new_n199_), .O(new_n596_));
  OR       g0580(.a(new_n596_), .b(i_2_5_91_0), .O(new_n597_));
  NAND     g0581(.a(new_n597_), .b(new_n170_), .O(new_n598_));
  OR       g0582(.a(new_n598_), .b(new_n595_), .O(new_n599_));
  OR       g0583(.a(new_n599_), .b(new_n593_), .O(new_n600_));
  AND      g0584(.a(new_n600_), .b(new_n20_), .O(new_n601_));
  OR       g0585(.a(new_n199_), .b(i_2_5_65_0), .O(new_n602_));
  NAND     g0586(.a(new_n602_), .b(new_n62_), .O(new_n603_));
  AND      g0587(.a(new_n190_), .b(i_2_5_102_0), .O(new_n604_));
  AND      g0588(.a(new_n604_), .b(new_n603_), .O(new_n605_));
  OR       g0589(.a(new_n178_), .b(i_2_5_148_0), .O(new_n606_));
  AND      g0590(.a(new_n352_), .b(new_n74_), .O(new_n607_));
  AND      g0591(.a(new_n607_), .b(new_n606_), .O(new_n608_));
  OR       g0592(.a(new_n608_), .b(new_n341_), .O(new_n609_));
  OR       g0593(.a(new_n609_), .b(new_n605_), .O(new_n610_));
  AND      g0594(.a(new_n610_), .b(new_n54_), .O(new_n611_));
  OR       g0595(.a(i_2_5_102_0), .b(new_n54_), .O(new_n612_));
  OR       g0596(.a(new_n276_), .b(new_n45_), .O(new_n613_));
  OR       g0597(.a(new_n613_), .b(new_n104_), .O(new_n614_));
  AND      g0598(.a(new_n614_), .b(new_n612_), .O(new_n615_));
  OR       g0599(.a(new_n295_), .b(new_n45_), .O(new_n616_));
  AND      g0600(.a(new_n616_), .b(i_2_5_82_0), .O(new_n617_));
  OR       g0601(.a(new_n563_), .b(new_n198_), .O(new_n618_));
  AND      g0602(.a(new_n618_), .b(new_n411_), .O(new_n619_));
  OR       g0603(.a(new_n619_), .b(new_n617_), .O(new_n620_));
  OR       g0604(.a(new_n620_), .b(new_n615_), .O(new_n621_));
  AND      g0605(.a(new_n621_), .b(i_2_5_12_0), .O(new_n622_));
  AND      g0606(.a(new_n176_), .b(i_2_5_148_0), .O(new_n623_));
  AND      g0607(.a(i_2_5_148_0), .b(new_n99_), .O(new_n624_));
  OR       g0608(.a(new_n624_), .b(new_n175_), .O(new_n625_));
  AND      g0609(.a(new_n625_), .b(new_n78_), .O(new_n626_));
  AND      g0610(.a(new_n626_), .b(new_n623_), .O(new_n627_));
  OR       g0611(.a(new_n627_), .b(new_n622_), .O(new_n628_));
  OR       g0612(.a(new_n628_), .b(new_n611_), .O(new_n629_));
  OR       g0613(.a(new_n629_), .b(new_n601_), .O(new_n630_));
  AND      g0614(.a(new_n630_), .b(new_n67_), .O(new_n631_));
  OR       g0615(.a(new_n326_), .b(new_n130_), .O(new_n632_));
  NAND     g0616(.a(new_n632_), .b(new_n602_), .O(new_n633_));
  OR       g0617(.a(new_n633_), .b(new_n499_), .O(new_n634_));
  AND      g0618(.a(new_n634_), .b(new_n72_), .O(new_n635_));
  OR       g0619(.a(new_n476_), .b(new_n65_), .O(new_n636_));
  AND      g0620(.a(new_n381_), .b(i_2_5_12_0), .O(new_n637_));
  NAND     g0621(.a(new_n637_), .b(new_n74_), .O(new_n638_));
  OR       g0622(.a(new_n638_), .b(new_n596_), .O(new_n639_));
  NAND     g0623(.a(new_n639_), .b(new_n636_), .O(new_n640_));
  OR       g0624(.a(new_n640_), .b(new_n635_), .O(new_n641_));
  AND      g0625(.a(new_n641_), .b(new_n54_), .O(new_n642_));
  AND      g0626(.a(new_n340_), .b(new_n51_), .O(new_n643_));
  NAND     g0627(.a(i_2_5_148_0), .b(i_2_5_12_0), .O(new_n644_));
  NOT      g0628(.a(new_n644_), .O(new_n645_));
  OR       g0629(.a(i_2_5_99_0), .b(i_2_5_82_0), .O(new_n646_));
  NAND     g0630(.a(new_n646_), .b(new_n113_), .O(new_n647_));
  AND      g0631(.a(new_n647_), .b(new_n645_), .O(new_n648_));
  OR       g0632(.a(new_n648_), .b(new_n643_), .O(new_n649_));
  OR       g0633(.a(new_n649_), .b(new_n642_), .O(new_n650_));
  AND      g0634(.a(new_n650_), .b(i_2_5_62_0), .O(new_n651_));
  NAND     g0635(.a(i_2_5_91_0), .b(i_2_5_70_0), .O(new_n652_));
  NOT      g0636(.a(new_n328_), .O(new_n653_));
  OR       g0637(.a(new_n499_), .b(i_2_5_12_0), .O(new_n654_));
  AND      g0638(.a(new_n654_), .b(new_n653_), .O(new_n655_));
  AND      g0639(.a(new_n364_), .b(new_n175_), .O(new_n656_));
  OR       g0640(.a(new_n656_), .b(new_n655_), .O(new_n657_));
  AND      g0641(.a(new_n657_), .b(new_n27_), .O(new_n658_));
  NAND     g0642(.a(new_n224_), .b(i_2_5_84_0), .O(new_n659_));
  NAND     g0643(.a(new_n659_), .b(new_n327_), .O(new_n660_));
  AND      g0644(.a(new_n660_), .b(new_n28_), .O(new_n661_));
  OR       g0645(.a(new_n661_), .b(new_n658_), .O(new_n662_));
  AND      g0646(.a(new_n662_), .b(new_n652_), .O(new_n663_));
  AND      g0647(.a(new_n652_), .b(new_n457_), .O(new_n664_));
  OR       g0648(.a(new_n328_), .b(new_n234_), .O(new_n665_));
  NOT      g0649(.a(new_n389_), .O(new_n666_));
  OR       g0650(.a(new_n666_), .b(new_n200_), .O(new_n667_));
  NAND     g0651(.a(new_n667_), .b(new_n665_), .O(new_n668_));
  OR       g0652(.a(new_n668_), .b(new_n664_), .O(new_n669_));
  AND      g0653(.a(new_n669_), .b(i_2_5_84_0), .O(new_n670_));
  AND      g0654(.a(new_n275_), .b(new_n54_), .O(new_n671_));
  AND      g0655(.a(i_2_5_82_0), .b(i_2_5_62_0), .O(new_n672_));
  OR       g0656(.a(new_n672_), .b(new_n45_), .O(new_n673_));
  AND      g0657(.a(i_2_5_148_0), .b(new_n67_), .O(new_n674_));
  AND      g0658(.a(new_n674_), .b(new_n673_), .O(new_n675_));
  OR       g0659(.a(new_n675_), .b(new_n160_), .O(new_n676_));
  AND      g0660(.a(new_n676_), .b(new_n345_), .O(new_n677_));
  OR       g0661(.a(new_n677_), .b(new_n671_), .O(new_n678_));
  OR       g0662(.a(new_n678_), .b(new_n670_), .O(new_n679_));
  OR       g0663(.a(new_n679_), .b(new_n663_), .O(new_n680_));
  OR       g0664(.a(new_n680_), .b(new_n651_), .O(new_n681_));
  OR       g0665(.a(new_n681_), .b(new_n631_), .O(new_n682_));
  OR       g0666(.a(new_n682_), .b(new_n590_), .O(new_n683_));
  AND      g0667(.a(new_n683_), .b(new_n21_), .O(new_n684_));
  NOT      g0668(.a(new_n602_), .O(new_n685_));
  OR       g0669(.a(i_2_5_102_0), .b(i_2_5_70_0), .O(new_n686_));
  AND      g0670(.a(new_n686_), .b(new_n685_), .O(new_n687_));
  OR       g0671(.a(new_n563_), .b(new_n295_), .O(new_n688_));
  AND      g0672(.a(new_n688_), .b(i_2_5_42_0), .O(new_n689_));
  OR       g0673(.a(new_n411_), .b(new_n51_), .O(new_n690_));
  AND      g0674(.a(new_n690_), .b(i_2_5_62_0), .O(new_n691_));
  OR       g0675(.a(new_n691_), .b(new_n689_), .O(new_n692_));
  AND      g0676(.a(new_n692_), .b(i_2_5_82_0), .O(new_n693_));
  OR       g0677(.a(new_n693_), .b(new_n687_), .O(new_n694_));
  AND      g0678(.a(new_n694_), .b(i_2_5_12_0), .O(new_n695_));
  AND      g0679(.a(new_n148_), .b(new_n27_), .O(new_n696_));
  OR       g0680(.a(new_n696_), .b(new_n660_), .O(new_n697_));
  AND      g0681(.a(new_n697_), .b(i_2_5_12_0), .O(new_n698_));
  OR       g0682(.a(new_n171_), .b(new_n118_), .O(new_n699_));
  AND      g0683(.a(new_n699_), .b(new_n623_), .O(new_n700_));
  OR       g0684(.a(new_n700_), .b(new_n300_), .O(new_n701_));
  OR       g0685(.a(new_n701_), .b(new_n698_), .O(new_n702_));
  AND      g0686(.a(new_n702_), .b(new_n54_), .O(new_n703_));
  AND      g0687(.a(new_n297_), .b(i_2_5_84_0), .O(new_n704_));
  AND      g0688(.a(new_n100_), .b(new_n54_), .O(new_n705_));
  OR       g0689(.a(new_n705_), .b(new_n704_), .O(new_n706_));
  AND      g0690(.a(new_n706_), .b(i_2_5_102_0), .O(new_n707_));
  OR       g0691(.a(new_n351_), .b(new_n313_), .O(new_n708_));
  AND      g0692(.a(new_n708_), .b(i_2_5_62_0), .O(new_n709_));
  OR       g0693(.a(new_n709_), .b(new_n216_), .O(new_n710_));
  OR       g0694(.a(new_n710_), .b(new_n707_), .O(new_n711_));
  AND      g0695(.a(new_n711_), .b(new_n450_), .O(new_n712_));
  AND      g0696(.a(new_n319_), .b(i_2_5_84_0), .O(new_n713_));
  AND      g0697(.a(new_n713_), .b(new_n563_), .O(new_n714_));
  OR       g0698(.a(new_n714_), .b(new_n712_), .O(new_n715_));
  OR       g0699(.a(new_n715_), .b(new_n703_), .O(new_n716_));
  OR       g0700(.a(new_n716_), .b(new_n695_), .O(new_n717_));
  AND      g0701(.a(new_n717_), .b(new_n20_), .O(new_n718_));
  AND      g0702(.a(new_n392_), .b(i_2_5_12_0), .O(new_n719_));
  AND      g0703(.a(new_n672_), .b(new_n34_), .O(new_n720_));
  OR       g0704(.a(new_n720_), .b(new_n719_), .O(new_n721_));
  AND      g0705(.a(new_n721_), .b(i_2_5_42_0), .O(new_n722_));
  AND      g0706(.a(new_n377_), .b(new_n27_), .O(new_n723_));
  AND      g0707(.a(new_n723_), .b(new_n215_), .O(new_n724_));
  OR       g0708(.a(new_n724_), .b(new_n722_), .O(new_n725_));
  AND      g0709(.a(new_n725_), .b(i_2_5_148_0), .O(new_n726_));
  OR       g0710(.a(new_n380_), .b(i_2_5_12_0), .O(new_n727_));
  AND      g0711(.a(new_n727_), .b(new_n79_), .O(new_n728_));
  OR       g0712(.a(new_n728_), .b(new_n726_), .O(new_n729_));
  AND      g0713(.a(new_n729_), .b(new_n55_), .O(new_n730_));
  OR       g0714(.a(new_n175_), .b(new_n54_), .O(new_n731_));
  NOT      g0715(.a(new_n131_), .O(new_n732_));
  NAND     g0716(.a(new_n602_), .b(i_2_5_70_0), .O(new_n733_));
  AND      g0717(.a(new_n733_), .b(new_n732_), .O(new_n734_));
  OR       g0718(.a(i_2_5_99_0), .b(i_2_5_70_0), .O(new_n735_));
  NOT      g0719(.a(new_n735_), .O(new_n736_));
  AND      g0720(.a(new_n736_), .b(i_2_5_148_0), .O(new_n737_));
  OR       g0721(.a(new_n737_), .b(new_n734_), .O(new_n738_));
  AND      g0722(.a(new_n738_), .b(i_2_5_82_0), .O(new_n739_));
  OR       g0723(.a(i_2_5_99_0), .b(new_n99_), .O(new_n740_));
  NOT      g0724(.a(new_n740_), .O(new_n741_));
  AND      g0725(.a(new_n741_), .b(new_n50_), .O(new_n742_));
  OR       g0726(.a(new_n742_), .b(new_n739_), .O(new_n743_));
  AND      g0727(.a(new_n743_), .b(new_n731_), .O(new_n744_));
  OR       g0728(.a(new_n72_), .b(i_2_5_82_0), .O(new_n745_));
  NOT      g0729(.a(new_n745_), .O(new_n746_));
  OR       g0730(.a(i_2_5_70_0), .b(i_2_5_65_0), .O(new_n747_));
  OR       g0731(.a(new_n747_), .b(new_n62_), .O(new_n748_));
  OR       g0732(.a(new_n748_), .b(new_n746_), .O(new_n749_));
  AND      g0733(.a(new_n749_), .b(new_n471_), .O(new_n750_));
  OR       g0734(.a(new_n750_), .b(new_n199_), .O(new_n751_));
  AND      g0735(.a(new_n118_), .b(new_n62_), .O(new_n752_));
  OR       g0736(.a(new_n518_), .b(new_n752_), .O(new_n753_));
  OR       g0737(.a(new_n753_), .b(new_n222_), .O(new_n754_));
  NAND     g0738(.a(new_n754_), .b(new_n751_), .O(new_n755_));
  AND      g0739(.a(new_n755_), .b(new_n86_), .O(new_n756_));
  OR       g0740(.a(new_n55_), .b(new_n20_), .O(new_n757_));
  OR       g0741(.a(new_n432_), .b(new_n261_), .O(new_n758_));
  NAND     g0742(.a(new_n758_), .b(new_n50_), .O(new_n759_));
  OR       g0743(.a(new_n753_), .b(new_n474_), .O(new_n760_));
  NAND     g0744(.a(new_n760_), .b(new_n759_), .O(new_n761_));
  AND      g0745(.a(new_n761_), .b(new_n757_), .O(new_n762_));
  OR       g0746(.a(new_n762_), .b(new_n756_), .O(new_n763_));
  OR       g0747(.a(new_n763_), .b(new_n744_), .O(new_n764_));
  OR       g0748(.a(new_n764_), .b(new_n730_), .O(new_n765_));
  OR       g0749(.a(new_n765_), .b(new_n718_), .O(new_n766_));
  OR       g0750(.a(new_n766_), .b(new_n684_), .O(new_n767_));
  OR       g0751(.a(new_n767_), .b(new_n514_), .O(new_n768_));
  OR       g0752(.a(new_n768_), .b(new_n274_), .O(new_n769_));
  AND      g0753(.a(new_n769_), .b(new_n18_), .O(new_n770_));
  AND      g0754(.a(new_n256_), .b(new_n19_), .O(new_n771_));
  OR       g0755(.a(new_n313_), .b(new_n55_), .O(new_n772_));
  AND      g0756(.a(new_n772_), .b(new_n190_), .O(new_n773_));
  NAND     g0757(.a(new_n740_), .b(new_n223_), .O(new_n774_));
  OR       g0758(.a(new_n774_), .b(new_n773_), .O(new_n775_));
  OR       g0759(.a(new_n775_), .b(new_n771_), .O(new_n776_));
  AND      g0760(.a(new_n776_), .b(i_2_5_84_0), .O(new_n777_));
  AND      g0761(.a(i_2_5_148_0), .b(i_2_5_42_0), .O(new_n778_));
  OR       g0762(.a(new_n778_), .b(new_n20_), .O(new_n779_));
  AND      g0763(.a(new_n779_), .b(new_n54_), .O(new_n780_));
  OR       g0764(.a(new_n780_), .b(new_n19_), .O(new_n781_));
  AND      g0765(.a(new_n297_), .b(i_2_5_102_0), .O(new_n782_));
  AND      g0766(.a(new_n782_), .b(new_n781_), .O(new_n783_));
  OR       g0767(.a(i_2_5_98_0), .b(i_2_5_65_0), .O(new_n784_));
  NOT      g0768(.a(new_n784_), .O(new_n785_));
  AND      g0769(.a(new_n54_), .b(i_2_5_12_0), .O(new_n786_));
  AND      g0770(.a(new_n786_), .b(i_2_5_84_0), .O(new_n787_));
  OR       g0771(.a(new_n787_), .b(new_n785_), .O(new_n788_));
  AND      g0772(.a(new_n788_), .b(new_n224_), .O(new_n789_));
  NOT      g0773(.a(new_n72_), .O(new_n790_));
  OR       g0774(.a(new_n602_), .b(new_n99_), .O(new_n791_));
  NAND     g0775(.a(new_n397_), .b(i_2_5_93_0), .O(new_n792_));
  NAND     g0776(.a(new_n792_), .b(new_n791_), .O(new_n793_));
  AND      g0777(.a(new_n793_), .b(new_n790_), .O(new_n794_));
  NAND     g0778(.a(new_n786_), .b(new_n563_), .O(new_n795_));
  OR       g0779(.a(i_2_5_98_0), .b(new_n130_), .O(new_n796_));
  OR       g0780(.a(new_n796_), .b(i_2_5_99_0), .O(new_n797_));
  NAND     g0781(.a(new_n797_), .b(new_n795_), .O(new_n798_));
  OR       g0782(.a(new_n798_), .b(new_n794_), .O(new_n799_));
  OR       g0783(.a(new_n799_), .b(new_n789_), .O(new_n800_));
  OR       g0784(.a(new_n800_), .b(new_n783_), .O(new_n801_));
  OR       g0785(.a(new_n801_), .b(new_n777_), .O(new_n802_));
  AND      g0786(.a(new_n802_), .b(i_2_5_82_0), .O(new_n803_));
  NAND     g0787(.a(new_n114_), .b(new_n199_), .O(new_n804_));
  OR       g0788(.a(new_n444_), .b(new_n20_), .O(new_n805_));
  OR       g0789(.a(new_n805_), .b(new_n448_), .O(new_n806_));
  AND      g0790(.a(new_n806_), .b(new_n804_), .O(new_n807_));
  OR       g0791(.a(new_n807_), .b(new_n298_), .O(new_n808_));
  AND      g0792(.a(new_n808_), .b(new_n19_), .O(new_n809_));
  OR       g0793(.a(i_2_5_99_0), .b(i_2_5_98_0), .O(new_n810_));
  NAND     g0794(.a(new_n810_), .b(new_n602_), .O(new_n811_));
  AND      g0795(.a(new_n811_), .b(new_n54_), .O(new_n812_));
  OR       g0796(.a(new_n812_), .b(new_n499_), .O(new_n813_));
  AND      g0797(.a(new_n813_), .b(new_n31_), .O(new_n814_));
  OR       g0798(.a(new_n65_), .b(i_2_5_98_0), .O(new_n815_));
  OR       g0799(.a(new_n815_), .b(new_n529_), .O(new_n816_));
  OR       g0800(.a(i_2_5_102_0), .b(new_n19_), .O(new_n817_));
  NAND     g0801(.a(new_n210_), .b(i_2_5_84_0), .O(new_n818_));
  OR       g0802(.a(new_n818_), .b(new_n817_), .O(new_n819_));
  NAND     g0803(.a(new_n819_), .b(new_n816_), .O(new_n820_));
  AND      g0804(.a(new_n820_), .b(new_n130_), .O(new_n821_));
  OR       g0805(.a(new_n113_), .b(new_n199_), .O(new_n822_));
  OR       g0806(.a(new_n646_), .b(new_n18_), .O(new_n823_));
  NAND     g0807(.a(new_n823_), .b(new_n822_), .O(new_n824_));
  AND      g0808(.a(new_n824_), .b(new_n426_), .O(new_n825_));
  OR       g0809(.a(new_n825_), .b(new_n821_), .O(new_n826_));
  OR       g0810(.a(new_n826_), .b(new_n814_), .O(new_n827_));
  OR       g0811(.a(new_n827_), .b(new_n809_), .O(new_n828_));
  OR       g0812(.a(new_n828_), .b(new_n803_), .O(new_n829_));
  AND      g0813(.a(new_n829_), .b(new_n21_), .O(new_n830_));
  AND      g0814(.a(new_n194_), .b(i_2_5_42_0), .O(new_n831_));
  NAND     g0815(.a(new_n381_), .b(new_n20_), .O(new_n832_));
  NAND     g0816(.a(new_n832_), .b(new_n815_), .O(new_n833_));
  OR       g0817(.a(new_n833_), .b(new_n831_), .O(new_n834_));
  AND      g0818(.a(new_n834_), .b(new_n27_), .O(new_n835_));
  NAND     g0819(.a(new_n644_), .b(i_2_5_99_0), .O(new_n836_));
  AND      g0820(.a(new_n836_), .b(i_2_5_84_0), .O(new_n837_));
  AND      g0821(.a(i_2_5_148_0), .b(new_n19_), .O(new_n838_));
  OR       g0822(.a(new_n838_), .b(new_n499_), .O(new_n839_));
  OR       g0823(.a(new_n839_), .b(new_n837_), .O(new_n840_));
  AND      g0824(.a(new_n840_), .b(i_2_5_102_0), .O(new_n841_));
  OR       g0825(.a(new_n444_), .b(new_n367_), .O(new_n842_));
  AND      g0826(.a(new_n842_), .b(new_n27_), .O(new_n843_));
  NAND     g0827(.a(new_n778_), .b(i_2_5_84_0), .O(new_n844_));
  OR       g0828(.a(new_n810_), .b(new_n99_), .O(new_n845_));
  NAND     g0829(.a(new_n845_), .b(new_n844_), .O(new_n846_));
  OR       g0830(.a(new_n846_), .b(new_n843_), .O(new_n847_));
  OR       g0831(.a(new_n847_), .b(new_n841_), .O(new_n848_));
  AND      g0832(.a(new_n848_), .b(new_n817_), .O(new_n849_));
  OR       g0833(.a(new_n849_), .b(new_n835_), .O(new_n850_));
  AND      g0834(.a(new_n850_), .b(new_n21_), .O(new_n851_));
  OR       g0835(.a(new_n51_), .b(i_2_5_12_0), .O(new_n852_));
  AND      g0836(.a(new_n852_), .b(new_n106_), .O(new_n853_));
  OR       g0837(.a(new_n853_), .b(new_n447_), .O(new_n854_));
  AND      g0838(.a(new_n854_), .b(i_2_5_102_0), .O(new_n855_));
  AND      g0839(.a(new_n282_), .b(new_n51_), .O(new_n856_));
  OR       g0840(.a(new_n458_), .b(new_n104_), .O(new_n857_));
  AND      g0841(.a(new_n857_), .b(new_n352_), .O(new_n858_));
  OR       g0842(.a(new_n858_), .b(new_n741_), .O(new_n859_));
  OR       g0843(.a(new_n859_), .b(new_n856_), .O(new_n860_));
  OR       g0844(.a(new_n860_), .b(new_n855_), .O(new_n861_));
  AND      g0845(.a(new_n861_), .b(i_2_5_148_0), .O(new_n862_));
  AND      g0846(.a(new_n280_), .b(new_n27_), .O(new_n863_));
  AND      g0847(.a(new_n20_), .b(i_2_5_84_0), .O(new_n864_));
  OR       g0848(.a(new_n864_), .b(i_2_5_12_0), .O(new_n865_));
  OR       g0849(.a(new_n865_), .b(new_n863_), .O(new_n866_));
  AND      g0850(.a(new_n106_), .b(i_2_5_102_0), .O(new_n867_));
  NAND     g0851(.a(new_n867_), .b(new_n866_), .O(new_n868_));
  NAND     g0852(.a(new_n868_), .b(new_n114_), .O(new_n869_));
  AND      g0853(.a(new_n869_), .b(i_2_5_82_0), .O(new_n870_));
  NAND     g0854(.a(i_2_5_98_0), .b(i_2_5_84_0), .O(new_n871_));
  OR       g0855(.a(new_n871_), .b(new_n186_), .O(new_n872_));
  NAND     g0856(.a(new_n872_), .b(new_n222_), .O(new_n873_));
  AND      g0857(.a(new_n873_), .b(new_n741_), .O(new_n874_));
  OR       g0858(.a(new_n874_), .b(new_n870_), .O(new_n875_));
  OR       g0859(.a(new_n875_), .b(new_n862_), .O(new_n876_));
  OR       g0860(.a(new_n876_), .b(new_n851_), .O(new_n877_));
  AND      g0861(.a(new_n877_), .b(new_n54_), .O(new_n878_));
  AND      g0862(.a(new_n745_), .b(new_n54_), .O(new_n879_));
  AND      g0863(.a(new_n75_), .b(i_2_5_82_0), .O(new_n880_));
  OR       g0864(.a(new_n880_), .b(new_n685_), .O(new_n881_));
  OR       g0865(.a(new_n881_), .b(new_n879_), .O(new_n882_));
  AND      g0866(.a(new_n882_), .b(i_2_5_12_0), .O(new_n883_));
  OR       g0867(.a(new_n563_), .b(new_n75_), .O(new_n884_));
  OR       g0868(.a(new_n884_), .b(new_n567_), .O(new_n885_));
  AND      g0869(.a(new_n885_), .b(new_n54_), .O(new_n886_));
  OR       g0870(.a(new_n27_), .b(i_2_5_42_0), .O(new_n887_));
  OR       g0871(.a(new_n276_), .b(new_n55_), .O(new_n888_));
  OR       g0872(.a(new_n888_), .b(new_n300_), .O(new_n889_));
  AND      g0873(.a(new_n889_), .b(new_n887_), .O(new_n890_));
  OR       g0874(.a(i_2_5_42_0), .b(i_2_5_12_0), .O(new_n891_));
  AND      g0875(.a(new_n891_), .b(new_n27_), .O(new_n892_));
  OR       g0876(.a(new_n892_), .b(i_2_5_148_0), .O(new_n893_));
  AND      g0877(.a(new_n612_), .b(new_n34_), .O(new_n894_));
  AND      g0878(.a(new_n894_), .b(new_n893_), .O(new_n895_));
  OR       g0879(.a(new_n895_), .b(new_n890_), .O(new_n896_));
  OR       g0880(.a(new_n896_), .b(new_n886_), .O(new_n897_));
  OR       g0881(.a(new_n897_), .b(new_n883_), .O(new_n898_));
  AND      g0882(.a(new_n898_), .b(new_n20_), .O(new_n899_));
  NOT      g0883(.a(new_n458_), .O(new_n900_));
  OR       g0884(.a(new_n568_), .b(new_n900_), .O(new_n901_));
  NAND     g0885(.a(i_2_5_93_0), .b(i_2_5_82_0), .O(new_n902_));
  OR       g0886(.a(new_n902_), .b(new_n530_), .O(new_n903_));
  NAND     g0887(.a(new_n903_), .b(new_n901_), .O(new_n904_));
  AND      g0888(.a(new_n904_), .b(new_n199_), .O(new_n905_));
  AND      g0889(.a(new_n891_), .b(new_n129_), .O(new_n906_));
  OR       g0890(.a(new_n906_), .b(new_n880_), .O(new_n907_));
  AND      g0891(.a(new_n907_), .b(new_n216_), .O(new_n908_));
  NAND     g0892(.a(new_n297_), .b(i_2_5_42_0), .O(new_n909_));
  NAND     g0893(.a(new_n909_), .b(new_n520_), .O(new_n910_));
  AND      g0894(.a(new_n910_), .b(new_n78_), .O(new_n911_));
  OR       g0895(.a(new_n911_), .b(new_n908_), .O(new_n912_));
  OR       g0896(.a(new_n912_), .b(new_n905_), .O(new_n913_));
  OR       g0897(.a(new_n913_), .b(new_n899_), .O(new_n914_));
  AND      g0898(.a(new_n914_), .b(new_n19_), .O(new_n915_));
  OR       g0899(.a(new_n170_), .b(new_n130_), .O(new_n916_));
  NAND     g0900(.a(new_n916_), .b(new_n900_), .O(new_n917_));
  OR       g0901(.a(i_2_5_82_0), .b(i_2_5_65_0), .O(new_n918_));
  AND      g0902(.a(new_n74_), .b(i_2_5_42_0), .O(new_n919_));
  AND      g0903(.a(new_n919_), .b(new_n918_), .O(new_n920_));
  OR       g0904(.a(new_n920_), .b(new_n52_), .O(new_n921_));
  AND      g0905(.a(new_n921_), .b(i_2_5_148_0), .O(new_n922_));
  OR       g0906(.a(new_n922_), .b(new_n917_), .O(new_n923_));
  AND      g0907(.a(new_n534_), .b(new_n191_), .O(new_n924_));
  AND      g0908(.a(new_n924_), .b(new_n923_), .O(new_n925_));
  AND      g0909(.a(new_n714_), .b(i_2_5_12_0), .O(new_n926_));
  OR       g0910(.a(new_n926_), .b(new_n925_), .O(new_n927_));
  OR       g0911(.a(new_n927_), .b(new_n915_), .O(new_n928_));
  OR       g0912(.a(new_n928_), .b(new_n878_), .O(new_n929_));
  OR       g0913(.a(new_n929_), .b(new_n830_), .O(new_n930_));
  AND      g0914(.a(new_n930_), .b(i_2_5_62_0), .O(new_n931_));
  OR       g0915(.a(new_n444_), .b(new_n423_), .O(new_n932_));
  AND      g0916(.a(new_n932_), .b(new_n21_), .O(new_n933_));
  OR       g0917(.a(new_n933_), .b(new_n58_), .O(new_n934_));
  AND      g0918(.a(new_n934_), .b(i_2_5_148_0), .O(new_n935_));
  OR       g0919(.a(i_2_5_148_0), .b(i_2_5_12_0), .O(new_n936_));
  NAND     g0920(.a(new_n936_), .b(new_n104_), .O(new_n937_));
  NOT      g0921(.a(new_n224_), .O(new_n938_));
  AND      g0922(.a(new_n407_), .b(new_n938_), .O(new_n939_));
  OR       g0923(.a(i_2_5_90_0), .b(new_n130_), .O(new_n940_));
  AND      g0924(.a(new_n940_), .b(i_2_5_99_0), .O(new_n941_));
  OR       g0925(.a(new_n229_), .b(new_n941_), .O(new_n942_));
  OR       g0926(.a(new_n942_), .b(new_n939_), .O(new_n943_));
  NAND     g0927(.a(new_n943_), .b(new_n937_), .O(new_n944_));
  OR       g0928(.a(new_n944_), .b(new_n935_), .O(new_n945_));
  AND      g0929(.a(new_n945_), .b(i_2_5_42_0), .O(new_n946_));
  AND      g0930(.a(i_2_5_148_0), .b(new_n21_), .O(new_n947_));
  OR       g0931(.a(new_n947_), .b(new_n20_), .O(new_n948_));
  AND      g0932(.a(new_n948_), .b(new_n171_), .O(new_n949_));
  OR       g0933(.a(new_n124_), .b(new_n104_), .O(new_n950_));
  AND      g0934(.a(new_n950_), .b(i_2_5_148_0), .O(new_n951_));
  OR       g0935(.a(new_n653_), .b(new_n124_), .O(new_n952_));
  AND      g0936(.a(new_n952_), .b(new_n21_), .O(new_n953_));
  OR       g0937(.a(new_n953_), .b(new_n951_), .O(new_n954_));
  AND      g0938(.a(new_n954_), .b(i_2_5_12_0), .O(new_n955_));
  OR       g0939(.a(new_n955_), .b(new_n949_), .O(new_n956_));
  OR       g0940(.a(new_n956_), .b(new_n946_), .O(new_n957_));
  AND      g0941(.a(new_n957_), .b(new_n27_), .O(new_n958_));
  OR       g0942(.a(new_n778_), .b(new_n470_), .O(new_n959_));
  AND      g0943(.a(new_n959_), .b(new_n228_), .O(new_n960_));
  NAND     g0944(.a(new_n279_), .b(new_n199_), .O(new_n961_));
  AND      g0945(.a(new_n961_), .b(new_n169_), .O(new_n962_));
  OR       g0946(.a(new_n864_), .b(new_n563_), .O(new_n963_));
  AND      g0947(.a(new_n963_), .b(new_n21_), .O(new_n964_));
  OR       g0948(.a(new_n964_), .b(new_n962_), .O(new_n965_));
  OR       g0949(.a(new_n965_), .b(new_n960_), .O(new_n966_));
  AND      g0950(.a(new_n199_), .b(i_2_5_93_0), .O(new_n967_));
  OR       g0951(.a(new_n500_), .b(new_n56_), .O(new_n968_));
  NAND     g0952(.a(new_n458_), .b(new_n65_), .O(new_n969_));
  NAND     g0953(.a(new_n969_), .b(new_n968_), .O(new_n970_));
  AND      g0954(.a(new_n970_), .b(new_n967_), .O(new_n971_));
  AND      g0955(.a(new_n31_), .b(i_2_5_148_0), .O(new_n972_));
  OR       g0956(.a(new_n972_), .b(new_n741_), .O(new_n973_));
  AND      g0957(.a(new_n973_), .b(new_n186_), .O(new_n974_));
  OR       g0958(.a(new_n974_), .b(new_n971_), .O(new_n975_));
  OR       g0959(.a(new_n975_), .b(new_n966_), .O(new_n976_));
  AND      g0960(.a(new_n976_), .b(new_n27_), .O(new_n977_));
  AND      g0961(.a(new_n194_), .b(new_n99_), .O(new_n978_));
  AND      g0962(.a(new_n426_), .b(new_n112_), .O(new_n979_));
  OR       g0963(.a(new_n979_), .b(new_n978_), .O(new_n980_));
  AND      g0964(.a(new_n980_), .b(i_2_5_82_0), .O(new_n981_));
  OR       g0965(.a(new_n563_), .b(new_n323_), .O(new_n982_));
  AND      g0966(.a(new_n224_), .b(new_n20_), .O(new_n983_));
  AND      g0967(.a(new_n983_), .b(new_n982_), .O(new_n984_));
  OR       g0968(.a(new_n984_), .b(new_n981_), .O(new_n985_));
  AND      g0969(.a(new_n985_), .b(new_n21_), .O(new_n986_));
  AND      g0970(.a(new_n917_), .b(new_n557_), .O(new_n987_));
  AND      g0971(.a(new_n28_), .b(i_2_5_102_0), .O(new_n988_));
  AND      g0972(.a(new_n72_), .b(i_2_5_42_0), .O(new_n989_));
  OR       g0973(.a(new_n989_), .b(new_n466_), .O(new_n990_));
  AND      g0974(.a(new_n990_), .b(i_2_5_148_0), .O(new_n991_));
  OR       g0975(.a(new_n991_), .b(new_n988_), .O(new_n992_));
  AND      g0976(.a(new_n992_), .b(new_n20_), .O(new_n993_));
  OR       g0977(.a(new_n993_), .b(new_n987_), .O(new_n994_));
  OR       g0978(.a(new_n994_), .b(new_n986_), .O(new_n995_));
  OR       g0979(.a(new_n995_), .b(new_n977_), .O(new_n996_));
  AND      g0980(.a(new_n996_), .b(new_n19_), .O(new_n997_));
  OR       g0981(.a(i_2_5_98_0), .b(i_2_5_90_0), .O(new_n998_));
  NOT      g0982(.a(new_n998_), .O(new_n999_));
  OR       g0983(.a(new_n999_), .b(new_n287_), .O(new_n1000_));
  AND      g0984(.a(new_n1000_), .b(new_n470_), .O(new_n1001_));
  AND      g0985(.a(new_n19_), .b(i_2_5_84_0), .O(new_n1002_));
  OR       g0986(.a(new_n1002_), .b(new_n466_), .O(new_n1003_));
  AND      g0987(.a(new_n1003_), .b(new_n21_), .O(new_n1004_));
  OR       g0988(.a(new_n1002_), .b(new_n50_), .O(new_n1005_));
  AND      g0989(.a(new_n1005_), .b(i_2_5_102_0), .O(new_n1006_));
  OR       g0990(.a(new_n1006_), .b(new_n1004_), .O(new_n1007_));
  AND      g0991(.a(new_n1007_), .b(i_2_5_82_0), .O(new_n1008_));
  OR       g0992(.a(new_n1008_), .b(new_n1001_), .O(new_n1009_));
  AND      g0993(.a(new_n1009_), .b(new_n779_), .O(new_n1010_));
  AND      g0994(.a(new_n323_), .b(i_2_5_12_0), .O(new_n1011_));
  AND      g0995(.a(new_n31_), .b(i_2_5_82_0), .O(new_n1012_));
  OR       g0996(.a(new_n1012_), .b(new_n1011_), .O(new_n1013_));
  NAND     g0997(.a(new_n170_), .b(i_2_5_90_0), .O(new_n1014_));
  AND      g0998(.a(new_n1014_), .b(new_n989_), .O(new_n1015_));
  OR       g0999(.a(new_n1015_), .b(new_n1013_), .O(new_n1016_));
  NAND     g1000(.a(new_n1016_), .b(new_n20_), .O(new_n1017_));
  NOT      g1001(.a(new_n28_), .O(new_n1018_));
  OR       g1002(.a(new_n142_), .b(new_n1018_), .O(new_n1019_));
  NAND     g1003(.a(new_n1019_), .b(new_n1017_), .O(new_n1020_));
  AND      g1004(.a(new_n1020_), .b(i_2_5_148_0), .O(new_n1021_));
  AND      g1005(.a(new_n1011_), .b(new_n196_), .O(new_n1022_));
  OR       g1006(.a(new_n1022_), .b(new_n1021_), .O(new_n1023_));
  OR       g1007(.a(new_n1023_), .b(new_n1010_), .O(new_n1024_));
  OR       g1008(.a(new_n1024_), .b(new_n997_), .O(new_n1025_));
  OR       g1009(.a(new_n1025_), .b(new_n958_), .O(new_n1026_));
  AND      g1010(.a(new_n1026_), .b(new_n54_), .O(new_n1027_));
  OR       g1011(.a(new_n40_), .b(i_2_5_148_0), .O(new_n1028_));
  NAND     g1012(.a(new_n948_), .b(new_n654_), .O(new_n1029_));
  NAND     g1013(.a(new_n1029_), .b(new_n1028_), .O(new_n1030_));
  AND      g1014(.a(new_n1030_), .b(i_2_5_82_0), .O(new_n1031_));
  NAND     g1015(.a(i_2_5_99_0), .b(i_2_5_82_0), .O(new_n1032_));
  AND      g1016(.a(new_n1032_), .b(new_n999_), .O(new_n1033_));
  OR       g1017(.a(i_2_5_148_0), .b(new_n130_), .O(new_n1034_));
  OR       g1018(.a(new_n1034_), .b(i_2_5_90_0), .O(new_n1035_));
  NAND     g1019(.a(new_n1035_), .b(new_n810_), .O(new_n1036_));
  AND      g1020(.a(new_n1036_), .b(new_n27_), .O(new_n1037_));
  OR       g1021(.a(new_n1037_), .b(new_n1033_), .O(new_n1038_));
  OR       g1022(.a(new_n1038_), .b(new_n1031_), .O(new_n1039_));
  AND      g1023(.a(new_n1039_), .b(i_2_5_42_0), .O(new_n1040_));
  AND      g1024(.a(new_n149_), .b(new_n221_), .O(new_n1041_));
  AND      g1025(.a(new_n1041_), .b(new_n19_), .O(new_n1042_));
  OR       g1026(.a(new_n326_), .b(i_2_5_98_0), .O(new_n1043_));
  NAND     g1027(.a(new_n1043_), .b(i_2_5_90_0), .O(new_n1044_));
  AND      g1028(.a(new_n1044_), .b(i_2_5_12_0), .O(new_n1045_));
  AND      g1029(.a(new_n624_), .b(new_n221_), .O(new_n1046_));
  AND      g1030(.a(new_n1046_), .b(new_n27_), .O(new_n1047_));
  OR       g1031(.a(new_n1047_), .b(new_n947_), .O(new_n1048_));
  OR       g1032(.a(new_n1048_), .b(new_n1045_), .O(new_n1049_));
  AND      g1033(.a(new_n1049_), .b(new_n20_), .O(new_n1050_));
  OR       g1034(.a(new_n1050_), .b(new_n1042_), .O(new_n1051_));
  OR       g1035(.a(new_n1051_), .b(new_n1040_), .O(new_n1052_));
  AND      g1036(.a(new_n1052_), .b(i_2_5_84_0), .O(new_n1053_));
  AND      g1037(.a(new_n28_), .b(i_2_5_148_0), .O(new_n1054_));
  OR       g1038(.a(new_n1054_), .b(new_n298_), .O(new_n1055_));
  AND      g1039(.a(new_n1055_), .b(new_n999_), .O(new_n1056_));
  NAND     g1040(.a(new_n998_), .b(new_n221_), .O(new_n1057_));
  AND      g1041(.a(new_n1057_), .b(new_n27_), .O(new_n1058_));
  AND      g1042(.a(new_n19_), .b(i_2_5_42_0), .O(new_n1059_));
  OR       g1043(.a(new_n1059_), .b(new_n21_), .O(new_n1060_));
  AND      g1044(.a(new_n1060_), .b(new_n248_), .O(new_n1061_));
  AND      g1045(.a(new_n1061_), .b(new_n1058_), .O(new_n1062_));
  OR       g1046(.a(new_n319_), .b(new_n21_), .O(new_n1063_));
  OR       g1047(.a(new_n1063_), .b(new_n785_), .O(new_n1064_));
  NAND     g1048(.a(new_n784_), .b(new_n199_), .O(new_n1065_));
  AND      g1049(.a(new_n481_), .b(i_2_5_12_0), .O(new_n1066_));
  AND      g1050(.a(new_n1066_), .b(new_n1065_), .O(new_n1067_));
  AND      g1051(.a(new_n1067_), .b(new_n1064_), .O(new_n1068_));
  OR       g1052(.a(new_n1068_), .b(new_n1062_), .O(new_n1069_));
  AND      g1053(.a(new_n1069_), .b(new_n20_), .O(new_n1070_));
  OR       g1054(.a(new_n1070_), .b(new_n1056_), .O(new_n1071_));
  OR       g1055(.a(new_n1071_), .b(new_n1053_), .O(new_n1072_));
  AND      g1056(.a(new_n1072_), .b(i_2_5_102_0), .O(new_n1073_));
  AND      g1057(.a(new_n499_), .b(new_n149_), .O(new_n1074_));
  AND      g1058(.a(new_n1074_), .b(i_2_5_91_0), .O(new_n1075_));
  NAND     g1059(.a(new_n298_), .b(new_n199_), .O(new_n1076_));
  OR       g1060(.a(new_n550_), .b(new_n130_), .O(new_n1077_));
  AND      g1061(.a(new_n1077_), .b(new_n1076_), .O(new_n1078_));
  OR       g1062(.a(new_n1078_), .b(i_2_5_90_0), .O(new_n1079_));
  OR       g1063(.a(new_n1011_), .b(new_n51_), .O(new_n1080_));
  AND      g1064(.a(new_n961_), .b(new_n191_), .O(new_n1081_));
  NAND     g1065(.a(new_n1081_), .b(new_n1080_), .O(new_n1082_));
  NAND     g1066(.a(new_n1082_), .b(new_n1079_), .O(new_n1083_));
  AND      g1067(.a(new_n1083_), .b(i_2_5_82_0), .O(new_n1084_));
  AND      g1068(.a(new_n21_), .b(i_2_5_65_0), .O(new_n1085_));
  AND      g1069(.a(new_n1085_), .b(new_n465_), .O(new_n1086_));
  OR       g1070(.a(new_n1086_), .b(new_n1084_), .O(new_n1087_));
  AND      g1071(.a(new_n1087_), .b(new_n19_), .O(new_n1088_));
  OR       g1072(.a(new_n1088_), .b(new_n1075_), .O(new_n1089_));
  OR       g1073(.a(new_n1089_), .b(new_n1073_), .O(new_n1090_));
  OR       g1074(.a(new_n1090_), .b(new_n1027_), .O(new_n1091_));
  OR       g1075(.a(new_n1091_), .b(new_n931_), .O(new_n1092_));
  AND      g1076(.a(new_n1092_), .b(new_n67_), .O(new_n1093_));
  OR       g1077(.a(new_n279_), .b(i_2_5_90_0), .O(new_n1094_));
  OR       g1078(.a(new_n1013_), .b(new_n319_), .O(new_n1095_));
  NAND     g1079(.a(new_n1095_), .b(i_2_5_102_0), .O(new_n1096_));
  NAND     g1080(.a(new_n1096_), .b(new_n1094_), .O(new_n1097_));
  AND      g1081(.a(new_n1097_), .b(new_n54_), .O(new_n1098_));
  NOT      g1082(.a(new_n967_), .O(new_n1099_));
  OR       g1083(.a(new_n1094_), .b(new_n1099_), .O(new_n1100_));
  AND      g1084(.a(new_n790_), .b(i_2_5_70_0), .O(new_n1101_));
  NAND     g1085(.a(new_n1101_), .b(new_n275_), .O(new_n1102_));
  NAND     g1086(.a(new_n1102_), .b(new_n1100_), .O(new_n1103_));
  AND      g1087(.a(new_n1103_), .b(new_n130_), .O(new_n1104_));
  AND      g1088(.a(new_n498_), .b(new_n92_), .O(new_n1105_));
  AND      g1089(.a(new_n196_), .b(i_2_5_42_0), .O(new_n1106_));
  OR       g1090(.a(new_n1106_), .b(new_n1105_), .O(new_n1107_));
  AND      g1091(.a(new_n1107_), .b(i_2_5_93_0), .O(new_n1108_));
  AND      g1092(.a(new_n550_), .b(new_n21_), .O(new_n1109_));
  AND      g1093(.a(new_n1109_), .b(new_n1012_), .O(new_n1110_));
  OR       g1094(.a(new_n1110_), .b(new_n1108_), .O(new_n1111_));
  OR       g1095(.a(new_n1111_), .b(new_n1104_), .O(new_n1112_));
  OR       g1096(.a(new_n1112_), .b(new_n1098_), .O(new_n1113_));
  AND      g1097(.a(new_n186_), .b(new_n54_), .O(new_n1114_));
  OR       g1098(.a(new_n988_), .b(new_n458_), .O(new_n1115_));
  OR       g1099(.a(new_n1115_), .b(new_n1114_), .O(new_n1116_));
  AND      g1100(.a(new_n1116_), .b(i_2_5_84_0), .O(new_n1117_));
  AND      g1101(.a(new_n500_), .b(new_n55_), .O(new_n1118_));
  OR       g1102(.a(new_n713_), .b(new_n149_), .O(new_n1119_));
  AND      g1103(.a(new_n1119_), .b(new_n65_), .O(new_n1120_));
  OR       g1104(.a(new_n1120_), .b(new_n1118_), .O(new_n1121_));
  OR       g1105(.a(new_n1121_), .b(new_n1117_), .O(new_n1122_));
  AND      g1106(.a(new_n1122_), .b(new_n20_), .O(new_n1123_));
  OR       g1107(.a(new_n787_), .b(new_n547_), .O(new_n1124_));
  AND      g1108(.a(new_n988_), .b(new_n112_), .O(new_n1125_));
  AND      g1109(.a(new_n757_), .b(new_n21_), .O(new_n1126_));
  OR       g1110(.a(new_n1126_), .b(new_n1125_), .O(new_n1127_));
  OR       g1111(.a(new_n1127_), .b(new_n1124_), .O(new_n1128_));
  OR       g1112(.a(new_n141_), .b(i_2_5_102_0), .O(new_n1129_));
  NAND     g1113(.a(new_n1129_), .b(new_n66_), .O(new_n1130_));
  AND      g1114(.a(new_n1130_), .b(i_2_5_42_0), .O(new_n1131_));
  OR       g1115(.a(new_n488_), .b(new_n18_), .O(new_n1132_));
  NAND     g1116(.a(new_n1132_), .b(new_n916_), .O(new_n1133_));
  AND      g1117(.a(new_n1133_), .b(new_n221_), .O(new_n1134_));
  OR       g1118(.a(new_n1134_), .b(new_n1131_), .O(new_n1135_));
  OR       g1119(.a(new_n1135_), .b(new_n1128_), .O(new_n1136_));
  AND      g1120(.a(new_n1136_), .b(i_2_5_148_0), .O(new_n1137_));
  OR       g1121(.a(new_n1137_), .b(new_n1123_), .O(new_n1138_));
  OR       g1122(.a(new_n1138_), .b(new_n1113_), .O(new_n1139_));
  AND      g1123(.a(new_n1139_), .b(new_n27_), .O(new_n1140_));
  AND      g1124(.a(new_n248_), .b(new_n20_), .O(new_n1141_));
  OR       g1125(.a(new_n947_), .b(new_n397_), .O(new_n1142_));
  AND      g1126(.a(new_n1142_), .b(i_2_5_42_0), .O(new_n1143_));
  OR       g1127(.a(new_n1143_), .b(new_n1141_), .O(new_n1144_));
  AND      g1128(.a(new_n1144_), .b(i_2_5_82_0), .O(new_n1145_));
  OR       g1129(.a(new_n1145_), .b(new_n501_), .O(new_n1146_));
  AND      g1130(.a(new_n1146_), .b(new_n54_), .O(new_n1147_));
  OR       g1131(.a(new_n499_), .b(new_n125_), .O(new_n1148_));
  NAND     g1132(.a(new_n1148_), .b(new_n339_), .O(new_n1149_));
  OR       g1133(.a(new_n199_), .b(i_2_5_90_0), .O(new_n1150_));
  AND      g1134(.a(new_n1150_), .b(new_n221_), .O(new_n1151_));
  AND      g1135(.a(new_n1150_), .b(i_2_5_99_0), .O(new_n1152_));
  OR       g1136(.a(new_n1152_), .b(new_n99_), .O(new_n1153_));
  OR       g1137(.a(new_n1153_), .b(new_n1151_), .O(new_n1154_));
  NAND     g1138(.a(new_n1154_), .b(new_n1149_), .O(new_n1155_));
  AND      g1139(.a(new_n1155_), .b(new_n54_), .O(new_n1156_));
  AND      g1140(.a(new_n551_), .b(i_2_5_42_0), .O(new_n1157_));
  OR       g1141(.a(new_n1157_), .b(new_n28_), .O(new_n1158_));
  AND      g1142(.a(new_n1158_), .b(new_n1141_), .O(new_n1159_));
  OR       g1143(.a(new_n313_), .b(new_n21_), .O(new_n1160_));
  OR       g1144(.a(i_2_5_148_0), .b(i_2_5_90_0), .O(new_n1161_));
  AND      g1145(.a(new_n221_), .b(i_2_5_12_0), .O(new_n1162_));
  AND      g1146(.a(new_n1162_), .b(new_n1161_), .O(new_n1163_));
  AND      g1147(.a(new_n1163_), .b(new_n1160_), .O(new_n1164_));
  OR       g1148(.a(new_n1164_), .b(new_n1159_), .O(new_n1165_));
  OR       g1149(.a(new_n1165_), .b(new_n1156_), .O(new_n1166_));
  AND      g1150(.a(new_n1166_), .b(i_2_5_84_0), .O(new_n1167_));
  OR       g1151(.a(new_n1167_), .b(new_n1147_), .O(new_n1168_));
  AND      g1152(.a(new_n1168_), .b(i_2_5_102_0), .O(new_n1169_));
  AND      g1153(.a(new_n481_), .b(i_2_5_84_0), .O(new_n1170_));
  OR       g1154(.a(new_n1170_), .b(new_n778_), .O(new_n1171_));
  AND      g1155(.a(new_n1171_), .b(new_n21_), .O(new_n1172_));
  NAND     g1156(.a(new_n338_), .b(new_n130_), .O(new_n1173_));
  OR       g1157(.a(new_n972_), .b(new_n22_), .O(new_n1174_));
  AND      g1158(.a(new_n1174_), .b(new_n1173_), .O(new_n1175_));
  OR       g1159(.a(new_n1175_), .b(new_n1172_), .O(new_n1176_));
  AND      g1160(.a(new_n1176_), .b(new_n20_), .O(new_n1177_));
  AND      g1161(.a(new_n99_), .b(i_2_5_12_0), .O(new_n1178_));
  AND      g1162(.a(new_n33_), .b(i_2_5_148_0), .O(new_n1179_));
  AND      g1163(.a(new_n1179_), .b(new_n1178_), .O(new_n1180_));
  OR       g1164(.a(new_n1180_), .b(new_n1177_), .O(new_n1181_));
  AND      g1165(.a(new_n1181_), .b(new_n54_), .O(new_n1182_));
  OR       g1166(.a(new_n1182_), .b(new_n1074_), .O(new_n1183_));
  OR       g1167(.a(new_n1183_), .b(new_n1169_), .O(new_n1184_));
  OR       g1168(.a(new_n1184_), .b(new_n1140_), .O(new_n1185_));
  AND      g1169(.a(new_n1185_), .b(i_2_5_62_0), .O(new_n1186_));
  OR       g1170(.a(new_n1178_), .b(new_n466_), .O(new_n1187_));
  AND      g1171(.a(new_n1187_), .b(new_n351_), .O(new_n1188_));
  AND      g1172(.a(new_n1171_), .b(i_2_5_102_0), .O(new_n1189_));
  AND      g1173(.a(new_n1178_), .b(i_2_5_148_0), .O(new_n1190_));
  AND      g1174(.a(new_n124_), .b(i_2_5_148_0), .O(new_n1191_));
  OR       g1175(.a(new_n1191_), .b(new_n988_), .O(new_n1192_));
  OR       g1176(.a(new_n1192_), .b(new_n1190_), .O(new_n1193_));
  OR       g1177(.a(new_n1193_), .b(new_n1189_), .O(new_n1194_));
  AND      g1178(.a(new_n1194_), .b(new_n21_), .O(new_n1195_));
  OR       g1179(.a(new_n1195_), .b(new_n1188_), .O(new_n1196_));
  AND      g1180(.a(new_n1196_), .b(new_n54_), .O(new_n1197_));
  AND      g1181(.a(new_n1179_), .b(new_n435_), .O(new_n1198_));
  OR       g1182(.a(i_2_5_90_0), .b(i_2_5_42_0), .O(new_n1199_));
  NAND     g1183(.a(new_n1199_), .b(new_n56_), .O(new_n1200_));
  OR       g1184(.a(new_n1200_), .b(new_n504_), .O(new_n1201_));
  AND      g1185(.a(new_n1201_), .b(i_2_5_148_0), .O(new_n1202_));
  AND      g1186(.a(new_n389_), .b(new_n21_), .O(new_n1203_));
  OR       g1187(.a(new_n1178_), .b(i_2_5_82_0), .O(new_n1204_));
  OR       g1188(.a(new_n1204_), .b(new_n1203_), .O(new_n1205_));
  AND      g1189(.a(new_n1205_), .b(new_n54_), .O(new_n1206_));
  OR       g1190(.a(new_n1206_), .b(new_n1202_), .O(new_n1207_));
  AND      g1191(.a(new_n1207_), .b(i_2_5_84_0), .O(new_n1208_));
  AND      g1192(.a(i_2_5_102_0), .b(new_n21_), .O(new_n1209_));
  OR       g1193(.a(new_n1209_), .b(i_2_5_148_0), .O(new_n1210_));
  AND      g1194(.a(new_n1114_), .b(i_2_5_42_0), .O(new_n1211_));
  OR       g1195(.a(new_n1211_), .b(new_n786_), .O(new_n1212_));
  AND      g1196(.a(new_n1212_), .b(new_n1210_), .O(new_n1213_));
  AND      g1197(.a(new_n343_), .b(new_n28_), .O(new_n1214_));
  AND      g1198(.a(new_n1209_), .b(i_2_5_148_0), .O(new_n1215_));
  OR       g1199(.a(new_n1215_), .b(new_n1214_), .O(new_n1216_));
  OR       g1200(.a(new_n1216_), .b(new_n1213_), .O(new_n1217_));
  OR       g1201(.a(new_n1217_), .b(new_n1208_), .O(new_n1218_));
  AND      g1202(.a(new_n1218_), .b(new_n27_), .O(new_n1219_));
  OR       g1203(.a(new_n1219_), .b(new_n1198_), .O(new_n1220_));
  OR       g1204(.a(new_n1220_), .b(new_n1197_), .O(new_n1221_));
  AND      g1205(.a(new_n1221_), .b(new_n20_), .O(new_n1222_));
  OR       g1206(.a(new_n644_), .b(new_n68_), .O(new_n1223_));
  NAND     g1207(.a(new_n1223_), .b(new_n131_), .O(new_n1224_));
  AND      g1208(.a(new_n1224_), .b(new_n434_), .O(new_n1225_));
  OR       g1209(.a(new_n1034_), .b(new_n112_), .O(new_n1226_));
  NAND     g1210(.a(new_n1226_), .b(new_n222_), .O(new_n1227_));
  AND      g1211(.a(new_n1227_), .b(i_2_5_42_0), .O(new_n1228_));
  OR       g1212(.a(new_n602_), .b(i_2_5_102_0), .O(new_n1229_));
  NAND     g1213(.a(new_n1229_), .b(new_n916_), .O(new_n1230_));
  OR       g1214(.a(new_n1230_), .b(new_n53_), .O(new_n1231_));
  OR       g1215(.a(new_n1231_), .b(new_n1228_), .O(new_n1232_));
  AND      g1216(.a(new_n1232_), .b(i_2_5_82_0), .O(new_n1233_));
  NAND     g1217(.a(new_n279_), .b(i_2_5_65_0), .O(new_n1234_));
  AND      g1218(.a(new_n852_), .b(new_n563_), .O(new_n1235_));
  AND      g1219(.a(new_n1235_), .b(new_n1234_), .O(new_n1236_));
  AND      g1220(.a(new_n1236_), .b(new_n446_), .O(new_n1237_));
  OR       g1221(.a(new_n1237_), .b(new_n1233_), .O(new_n1238_));
  AND      g1222(.a(new_n1238_), .b(new_n21_), .O(new_n1239_));
  OR       g1223(.a(new_n1239_), .b(new_n1225_), .O(new_n1240_));
  AND      g1224(.a(new_n1240_), .b(new_n54_), .O(new_n1241_));
  NOT      g1225(.a(new_n142_), .O(new_n1242_));
  NOT      g1226(.a(new_n1032_), .O(new_n1243_));
  AND      g1227(.a(new_n1243_), .b(new_n458_), .O(new_n1244_));
  AND      g1228(.a(new_n1244_), .b(new_n1242_), .O(new_n1245_));
  OR       g1229(.a(new_n1245_), .b(new_n1241_), .O(new_n1246_));
  OR       g1230(.a(new_n1246_), .b(new_n1222_), .O(new_n1247_));
  OR       g1231(.a(new_n1247_), .b(new_n1186_), .O(new_n1248_));
  AND      g1232(.a(new_n1248_), .b(new_n19_), .O(new_n1249_));
  OR       g1233(.a(new_n351_), .b(new_n323_), .O(new_n1250_));
  NAND     g1234(.a(new_n338_), .b(i_2_5_90_0), .O(new_n1251_));
  AND      g1235(.a(new_n1251_), .b(i_2_5_62_0), .O(new_n1252_));
  AND      g1236(.a(new_n1252_), .b(new_n1250_), .O(new_n1253_));
  OR       g1237(.a(new_n1253_), .b(new_n1179_), .O(new_n1254_));
  AND      g1238(.a(new_n1254_), .b(new_n1170_), .O(new_n1255_));
  OR       g1239(.a(new_n1255_), .b(i_2_5_12_0), .O(new_n1256_));
  NOT      g1240(.a(new_n1170_), .O(new_n1257_));
  NAND     g1241(.a(new_n1257_), .b(new_n791_), .O(new_n1258_));
  OR       g1242(.a(new_n1258_), .b(new_n1253_), .O(new_n1259_));
  AND      g1243(.a(new_n1259_), .b(new_n1256_), .O(new_n1260_));
  OR       g1244(.a(new_n1041_), .b(new_n685_), .O(new_n1261_));
  AND      g1245(.a(new_n1261_), .b(new_n392_), .O(new_n1262_));
  NAND     g1246(.a(new_n1150_), .b(new_n566_), .O(new_n1263_));
  OR       g1247(.a(new_n1263_), .b(new_n1253_), .O(new_n1264_));
  AND      g1248(.a(new_n1264_), .b(new_n27_), .O(new_n1265_));
  OR       g1249(.a(new_n1265_), .b(new_n1262_), .O(new_n1266_));
  OR       g1250(.a(new_n1266_), .b(new_n1260_), .O(new_n1267_));
  AND      g1251(.a(new_n1267_), .b(i_2_5_102_0), .O(new_n1268_));
  AND      g1252(.a(new_n232_), .b(i_2_5_12_0), .O(new_n1269_));
  OR       g1253(.a(i_2_5_62_0), .b(i_2_5_42_0), .O(new_n1270_));
  AND      g1254(.a(new_n1270_), .b(new_n23_), .O(new_n1271_));
  OR       g1255(.a(new_n1271_), .b(new_n1269_), .O(new_n1272_));
  AND      g1256(.a(new_n1272_), .b(new_n27_), .O(new_n1273_));
  AND      g1257(.a(new_n352_), .b(new_n149_), .O(new_n1274_));
  OR       g1258(.a(new_n1274_), .b(new_n1273_), .O(new_n1275_));
  AND      g1259(.a(new_n1275_), .b(i_2_5_148_0), .O(new_n1276_));
  NAND     g1260(.a(new_n1179_), .b(new_n99_), .O(new_n1277_));
  NAND     g1261(.a(new_n1277_), .b(new_n144_), .O(new_n1278_));
  AND      g1262(.a(new_n1278_), .b(new_n72_), .O(new_n1279_));
  OR       g1263(.a(new_n465_), .b(new_n41_), .O(new_n1280_));
  AND      g1264(.a(new_n1280_), .b(new_n672_), .O(new_n1281_));
  OR       g1265(.a(new_n1281_), .b(new_n1279_), .O(new_n1282_));
  OR       g1266(.a(new_n1282_), .b(new_n1276_), .O(new_n1283_));
  OR       g1267(.a(new_n1283_), .b(new_n1268_), .O(new_n1284_));
  AND      g1268(.a(new_n1284_), .b(new_n54_), .O(new_n1285_));
  NAND     g1269(.a(i_2_5_93_0), .b(i_2_5_70_0), .O(new_n1286_));
  OR       g1270(.a(new_n1286_), .b(new_n1150_), .O(new_n1287_));
  NAND     g1271(.a(new_n300_), .b(i_2_5_98_0), .O(new_n1288_));
  NAND     g1272(.a(new_n1288_), .b(new_n1287_), .O(new_n1289_));
  AND      g1273(.a(new_n1289_), .b(i_2_5_42_0), .O(new_n1290_));
  AND      g1274(.a(i_2_5_98_0), .b(i_2_5_12_0), .O(new_n1291_));
  OR       g1275(.a(new_n1291_), .b(new_n21_), .O(new_n1292_));
  AND      g1276(.a(new_n1292_), .b(new_n563_), .O(new_n1293_));
  OR       g1277(.a(new_n1293_), .b(new_n1290_), .O(new_n1294_));
  AND      g1278(.a(new_n1294_), .b(new_n27_), .O(new_n1295_));
  AND      g1279(.a(new_n33_), .b(new_n65_), .O(new_n1296_));
  OR       g1280(.a(new_n1296_), .b(new_n563_), .O(new_n1297_));
  AND      g1281(.a(new_n112_), .b(i_2_5_42_0), .O(new_n1298_));
  AND      g1282(.a(new_n1298_), .b(new_n1297_), .O(new_n1299_));
  OR       g1283(.a(new_n1299_), .b(new_n1215_), .O(new_n1300_));
  AND      g1284(.a(new_n1300_), .b(i_2_5_12_0), .O(new_n1301_));
  AND      g1285(.a(i_2_5_98_0), .b(i_2_5_93_0), .O(new_n1302_));
  AND      g1286(.a(new_n1302_), .b(new_n426_), .O(new_n1303_));
  AND      g1287(.a(new_n1303_), .b(new_n947_), .O(new_n1304_));
  OR       g1288(.a(new_n1304_), .b(new_n1301_), .O(new_n1305_));
  OR       g1289(.a(new_n1305_), .b(new_n1295_), .O(new_n1306_));
  AND      g1290(.a(new_n1306_), .b(i_2_5_62_0), .O(new_n1307_));
  NAND     g1291(.a(new_n936_), .b(i_2_5_82_0), .O(new_n1308_));
  NAND     g1292(.a(new_n1308_), .b(new_n916_), .O(new_n1309_));
  AND      g1293(.a(new_n1309_), .b(new_n41_), .O(new_n1310_));
  OR       g1294(.a(new_n1310_), .b(new_n1307_), .O(new_n1311_));
  OR       g1295(.a(new_n1311_), .b(new_n1285_), .O(new_n1312_));
  AND      g1296(.a(new_n1312_), .b(new_n20_), .O(new_n1313_));
  AND      g1297(.a(new_n118_), .b(new_n22_), .O(new_n1314_));
  NOT      g1298(.a(new_n795_), .O(new_n1315_));
  AND      g1299(.a(new_n1315_), .b(i_2_5_62_0), .O(new_n1316_));
  AND      g1300(.a(new_n1316_), .b(new_n1314_), .O(new_n1317_));
  OR       g1301(.a(new_n423_), .b(new_n171_), .O(new_n1318_));
  AND      g1302(.a(new_n1318_), .b(new_n216_), .O(new_n1319_));
  AND      g1303(.a(i_2_5_99_0), .b(new_n221_), .O(new_n1320_));
  AND      g1304(.a(new_n786_), .b(new_n1320_), .O(new_n1321_));
  OR       g1305(.a(new_n1321_), .b(new_n1054_), .O(new_n1322_));
  OR       g1306(.a(new_n1322_), .b(new_n1319_), .O(new_n1323_));
  AND      g1307(.a(new_n1323_), .b(i_2_5_62_0), .O(new_n1324_));
  AND      g1308(.a(new_n972_), .b(new_n55_), .O(new_n1325_));
  AND      g1309(.a(new_n1325_), .b(new_n932_), .O(new_n1326_));
  OR       g1310(.a(new_n1326_), .b(new_n1324_), .O(new_n1327_));
  AND      g1311(.a(new_n1327_), .b(i_2_5_42_0), .O(new_n1328_));
  AND      g1312(.a(new_n262_), .b(new_n161_), .O(new_n1329_));
  AND      g1313(.a(new_n625_), .b(new_n28_), .O(new_n1330_));
  OR       g1314(.a(new_n1330_), .b(new_n1329_), .O(new_n1331_));
  AND      g1315(.a(new_n1331_), .b(new_n295_), .O(new_n1332_));
  OR       g1316(.a(new_n1332_), .b(new_n1328_), .O(new_n1333_));
  AND      g1317(.a(new_n1333_), .b(new_n21_), .O(new_n1334_));
  NOT      g1318(.a(new_n902_), .O(new_n1335_));
  OR       g1319(.a(new_n1335_), .b(new_n433_), .O(new_n1336_));
  AND      g1320(.a(new_n645_), .b(new_n122_), .O(new_n1337_));
  AND      g1321(.a(new_n1337_), .b(new_n1336_), .O(new_n1338_));
  OR       g1322(.a(new_n1338_), .b(new_n1334_), .O(new_n1339_));
  AND      g1323(.a(new_n1339_), .b(new_n27_), .O(new_n1340_));
  OR       g1324(.a(new_n1340_), .b(new_n1317_), .O(new_n1341_));
  OR       g1325(.a(new_n1341_), .b(new_n1313_), .O(new_n1342_));
  OR       g1326(.a(new_n1342_), .b(new_n1249_), .O(new_n1343_));
  OR       g1327(.a(new_n1343_), .b(new_n1093_), .O(new_n1344_));
  OR       g1328(.a(new_n1344_), .b(new_n770_), .O(new_n1345_));
  AND      g1329(.a(new_n1345_), .b(new_n17_), .O(new_n1346_));
  AND      g1330(.a(i_2_5_62_0), .b(new_n99_), .O(new_n1347_));
  AND      g1331(.a(new_n1347_), .b(i_2_5_98_0), .O(new_n1348_));
  OR       g1332(.a(new_n1348_), .b(new_n1059_), .O(new_n1349_));
  AND      g1333(.a(new_n1349_), .b(new_n130_), .O(new_n1350_));
  AND      g1334(.a(new_n19_), .b(i_2_5_12_0), .O(new_n1351_));
  OR       g1335(.a(new_n1351_), .b(new_n21_), .O(new_n1352_));
  AND      g1336(.a(new_n1352_), .b(i_2_5_62_0), .O(new_n1353_));
  OR       g1337(.a(new_n1353_), .b(new_n196_), .O(new_n1354_));
  OR       g1338(.a(new_n1354_), .b(new_n1350_), .O(new_n1355_));
  AND      g1339(.a(new_n1355_), .b(new_n67_), .O(new_n1356_));
  NAND     g1340(.a(new_n229_), .b(new_n180_), .O(new_n1357_));
  AND      g1341(.a(new_n1357_), .b(new_n19_), .O(new_n1358_));
  NOT      g1342(.a(new_n810_), .O(new_n1359_));
  AND      g1343(.a(new_n21_), .b(i_2_5_62_0), .O(new_n1360_));
  OR       g1344(.a(new_n1360_), .b(new_n1359_), .O(new_n1361_));
  AND      g1345(.a(new_n1361_), .b(i_2_5_12_0), .O(new_n1362_));
  OR       g1346(.a(new_n1362_), .b(new_n250_), .O(new_n1363_));
  OR       g1347(.a(new_n1363_), .b(new_n1358_), .O(new_n1364_));
  OR       g1348(.a(new_n1364_), .b(new_n1356_), .O(new_n1365_));
  AND      g1349(.a(new_n1365_), .b(i_2_5_148_0), .O(new_n1366_));
  OR       g1350(.a(new_n998_), .b(new_n67_), .O(new_n1367_));
  OR       g1351(.a(new_n1367_), .b(new_n31_), .O(new_n1368_));
  NAND     g1352(.a(new_n1368_), .b(new_n143_), .O(new_n1369_));
  AND      g1353(.a(new_n1369_), .b(i_2_5_82_0), .O(new_n1370_));
  AND      g1354(.a(new_n149_), .b(new_n67_), .O(new_n1371_));
  AND      g1355(.a(new_n19_), .b(i_2_5_62_0), .O(new_n1372_));
  OR       g1356(.a(new_n1372_), .b(new_n1351_), .O(new_n1373_));
  OR       g1357(.a(new_n1373_), .b(new_n1371_), .O(new_n1374_));
  NAND     g1358(.a(i_2_5_90_0), .b(i_2_5_70_0), .O(new_n1375_));
  AND      g1359(.a(new_n1375_), .b(new_n20_), .O(new_n1376_));
  AND      g1360(.a(new_n1376_), .b(new_n1374_), .O(new_n1377_));
  OR       g1361(.a(new_n1377_), .b(new_n1370_), .O(new_n1378_));
  AND      g1362(.a(new_n1378_), .b(i_2_5_42_0), .O(new_n1379_));
  AND      g1363(.a(new_n457_), .b(new_n29_), .O(new_n1380_));
  AND      g1364(.a(new_n19_), .b(i_2_5_82_0), .O(new_n1381_));
  OR       g1365(.a(new_n1381_), .b(i_2_5_12_0), .O(new_n1382_));
  AND      g1366(.a(i_2_5_99_0), .b(i_2_5_90_0), .O(new_n1383_));
  NOT      g1367(.a(new_n1383_), .O(new_n1384_));
  AND      g1368(.a(new_n1384_), .b(new_n1382_), .O(new_n1385_));
  AND      g1369(.a(new_n1291_), .b(new_n199_), .O(new_n1386_));
  OR       g1370(.a(new_n1386_), .b(new_n196_), .O(new_n1387_));
  OR       g1371(.a(new_n1387_), .b(new_n1385_), .O(new_n1388_));
  AND      g1372(.a(new_n1388_), .b(new_n67_), .O(new_n1389_));
  OR       g1373(.a(new_n1389_), .b(new_n1380_), .O(new_n1390_));
  AND      g1374(.a(new_n1390_), .b(i_2_5_62_0), .O(new_n1391_));
  OR       g1375(.a(i_2_5_90_0), .b(i_2_5_70_0), .O(new_n1392_));
  NOT      g1376(.a(new_n1392_), .O(new_n1393_));
  AND      g1377(.a(new_n112_), .b(i_2_5_62_0), .O(new_n1394_));
  AND      g1378(.a(new_n1394_), .b(new_n1393_), .O(new_n1395_));
  AND      g1379(.a(new_n1395_), .b(i_2_5_98_0), .O(new_n1396_));
  AND      g1380(.a(new_n19_), .b(i_2_5_90_0), .O(new_n1397_));
  AND      g1381(.a(new_n1397_), .b(new_n1190_), .O(new_n1398_));
  OR       g1382(.a(new_n1398_), .b(new_n1396_), .O(new_n1399_));
  AND      g1383(.a(new_n1399_), .b(new_n221_), .O(new_n1400_));
  OR       g1384(.a(new_n999_), .b(new_n28_), .O(new_n1401_));
  AND      g1385(.a(new_n1401_), .b(new_n736_), .O(new_n1402_));
  OR       g1386(.a(new_n1402_), .b(new_n1400_), .O(new_n1403_));
  OR       g1387(.a(new_n1403_), .b(new_n1391_), .O(new_n1404_));
  OR       g1388(.a(new_n1404_), .b(new_n1379_), .O(new_n1405_));
  OR       g1389(.a(new_n1405_), .b(new_n1366_), .O(new_n1406_));
  AND      g1390(.a(new_n1406_), .b(new_n27_), .O(new_n1407_));
  OR       g1391(.a(new_n534_), .b(new_n19_), .O(new_n1408_));
  OR       g1392(.a(new_n1408_), .b(new_n68_), .O(new_n1409_));
  OR       g1393(.a(new_n199_), .b(i_2_5_98_0), .O(new_n1410_));
  AND      g1394(.a(new_n1410_), .b(new_n526_), .O(new_n1411_));
  NAND     g1395(.a(new_n1411_), .b(new_n1409_), .O(new_n1412_));
  AND      g1396(.a(new_n1412_), .b(i_2_5_42_0), .O(new_n1413_));
  AND      g1397(.a(new_n190_), .b(new_n19_), .O(new_n1414_));
  AND      g1398(.a(new_n1414_), .b(new_n733_), .O(new_n1415_));
  OR       g1399(.a(new_n1415_), .b(new_n1413_), .O(new_n1416_));
  AND      g1400(.a(new_n1416_), .b(new_n21_), .O(new_n1417_));
  AND      g1401(.a(new_n1060_), .b(i_2_5_148_0), .O(new_n1418_));
  OR       g1402(.a(new_n21_), .b(i_2_5_82_0), .O(new_n1419_));
  OR       g1403(.a(i_2_5_98_0), .b(i_2_5_70_0), .O(new_n1420_));
  NOT      g1404(.a(new_n1420_), .O(new_n1421_));
  AND      g1405(.a(new_n1421_), .b(new_n1419_), .O(new_n1422_));
  OR       g1406(.a(new_n1422_), .b(new_n1418_), .O(new_n1423_));
  OR       g1407(.a(i_2_5_82_0), .b(i_2_5_70_0), .O(new_n1424_));
  NAND     g1408(.a(new_n1424_), .b(new_n998_), .O(new_n1425_));
  AND      g1409(.a(new_n1425_), .b(i_2_5_42_0), .O(new_n1426_));
  NAND     g1410(.a(new_n784_), .b(new_n130_), .O(new_n1427_));
  AND      g1411(.a(new_n1427_), .b(new_n1375_), .O(new_n1428_));
  OR       g1412(.a(new_n1059_), .b(i_2_5_82_0), .O(new_n1429_));
  AND      g1413(.a(new_n1429_), .b(new_n27_), .O(new_n1430_));
  OR       g1414(.a(new_n1430_), .b(new_n1428_), .O(new_n1431_));
  OR       g1415(.a(new_n1431_), .b(new_n1426_), .O(new_n1432_));
  OR       g1416(.a(new_n1432_), .b(new_n1423_), .O(new_n1433_));
  AND      g1417(.a(new_n1433_), .b(new_n20_), .O(new_n1434_));
  OR       g1418(.a(new_n1434_), .b(new_n1417_), .O(new_n1435_));
  AND      g1419(.a(new_n1435_), .b(i_2_5_62_0), .O(new_n1436_));
  OR       g1420(.a(new_n796_), .b(new_n20_), .O(new_n1437_));
  NAND     g1421(.a(new_n1437_), .b(new_n735_), .O(new_n1438_));
  AND      g1422(.a(new_n1438_), .b(new_n221_), .O(new_n1439_));
  AND      g1423(.a(new_n1065_), .b(new_n20_), .O(new_n1440_));
  OR       g1424(.a(new_n1440_), .b(new_n1439_), .O(new_n1441_));
  AND      g1425(.a(new_n1441_), .b(i_2_5_42_0), .O(new_n1442_));
  NAND     g1426(.a(new_n1420_), .b(i_2_5_65_0), .O(new_n1443_));
  AND      g1427(.a(new_n1443_), .b(new_n210_), .O(new_n1444_));
  OR       g1428(.a(new_n1381_), .b(i_2_5_148_0), .O(new_n1445_));
  AND      g1429(.a(new_n1445_), .b(new_n67_), .O(new_n1446_));
  AND      g1430(.a(new_n1381_), .b(new_n190_), .O(new_n1447_));
  OR       g1431(.a(new_n1447_), .b(new_n278_), .O(new_n1448_));
  OR       g1432(.a(new_n1448_), .b(new_n1446_), .O(new_n1449_));
  AND      g1433(.a(new_n1449_), .b(i_2_5_12_0), .O(new_n1450_));
  OR       g1434(.a(new_n1450_), .b(new_n1444_), .O(new_n1451_));
  OR       g1435(.a(new_n1451_), .b(new_n1442_), .O(new_n1452_));
  AND      g1436(.a(new_n1452_), .b(new_n21_), .O(new_n1453_));
  OR       g1437(.a(new_n602_), .b(new_n21_), .O(new_n1454_));
  OR       g1438(.a(new_n747_), .b(new_n99_), .O(new_n1455_));
  AND      g1439(.a(new_n1455_), .b(new_n797_), .O(new_n1456_));
  NAND     g1440(.a(new_n1456_), .b(new_n1454_), .O(new_n1457_));
  AND      g1441(.a(new_n1457_), .b(i_2_5_82_0), .O(new_n1458_));
  AND      g1442(.a(new_n654_), .b(i_2_5_42_0), .O(new_n1459_));
  OR       g1443(.a(i_2_5_65_0), .b(i_2_5_42_0), .O(new_n1460_));
  NAND     g1444(.a(new_n1460_), .b(new_n796_), .O(new_n1461_));
  AND      g1445(.a(new_n1461_), .b(i_2_5_148_0), .O(new_n1462_));
  OR       g1446(.a(new_n1462_), .b(new_n1459_), .O(new_n1463_));
  AND      g1447(.a(new_n1463_), .b(new_n67_), .O(new_n1464_));
  OR       g1448(.a(i_2_5_70_0), .b(i_2_5_62_0), .O(new_n1465_));
  NOT      g1449(.a(new_n1465_), .O(new_n1466_));
  OR       g1450(.a(new_n1466_), .b(new_n250_), .O(new_n1467_));
  AND      g1451(.a(new_n838_), .b(i_2_5_82_0), .O(new_n1468_));
  OR       g1452(.a(new_n1468_), .b(new_n50_), .O(new_n1469_));
  AND      g1453(.a(new_n1469_), .b(new_n1467_), .O(new_n1470_));
  AND      g1454(.a(new_n1360_), .b(new_n100_), .O(new_n1471_));
  OR       g1455(.a(new_n1471_), .b(new_n645_), .O(new_n1472_));
  AND      g1456(.a(new_n1472_), .b(new_n20_), .O(new_n1473_));
  OR       g1457(.a(new_n1473_), .b(new_n1470_), .O(new_n1474_));
  OR       g1458(.a(new_n1474_), .b(new_n1464_), .O(new_n1475_));
  OR       g1459(.a(new_n1475_), .b(new_n1458_), .O(new_n1476_));
  OR       g1460(.a(new_n1476_), .b(new_n1453_), .O(new_n1477_));
  OR       g1461(.a(new_n1477_), .b(new_n1436_), .O(new_n1478_));
  AND      g1462(.a(new_n1478_), .b(i_2_5_84_0), .O(new_n1479_));
  OR       g1463(.a(i_2_5_98_0), .b(new_n27_), .O(new_n1480_));
  OR       g1464(.a(new_n1480_), .b(new_n31_), .O(new_n1481_));
  NAND     g1465(.a(new_n1481_), .b(new_n551_), .O(new_n1482_));
  AND      g1466(.a(new_n1482_), .b(i_2_5_62_0), .O(new_n1483_));
  AND      g1467(.a(new_n112_), .b(i_2_5_82_0), .O(new_n1484_));
  OR       g1468(.a(new_n1484_), .b(new_n1351_), .O(new_n1485_));
  AND      g1469(.a(new_n1485_), .b(new_n20_), .O(new_n1486_));
  OR       g1470(.a(new_n1486_), .b(new_n1483_), .O(new_n1487_));
  AND      g1471(.a(new_n1487_), .b(i_2_5_42_0), .O(new_n1488_));
  OR       g1472(.a(new_n838_), .b(new_n250_), .O(new_n1489_));
  AND      g1473(.a(new_n1489_), .b(i_2_5_12_0), .O(new_n1490_));
  OR       g1474(.a(new_n1490_), .b(new_n1488_), .O(new_n1491_));
  AND      g1475(.a(new_n1491_), .b(new_n21_), .O(new_n1492_));
  OR       g1476(.a(i_2_5_98_0), .b(new_n221_), .O(new_n1493_));
  NAND     g1477(.a(new_n1493_), .b(new_n1034_), .O(new_n1494_));
  AND      g1478(.a(new_n1494_), .b(i_2_5_42_0), .O(new_n1495_));
  OR       g1479(.a(new_n1173_), .b(new_n999_), .O(new_n1496_));
  OR       g1480(.a(new_n1496_), .b(new_n1495_), .O(new_n1497_));
  OR       g1481(.a(new_n672_), .b(i_2_5_148_0), .O(new_n1498_));
  AND      g1482(.a(new_n1498_), .b(new_n20_), .O(new_n1499_));
  AND      g1483(.a(new_n1499_), .b(new_n1497_), .O(new_n1500_));
  OR       g1484(.a(new_n1500_), .b(new_n1492_), .O(new_n1501_));
  AND      g1485(.a(new_n1501_), .b(new_n67_), .O(new_n1502_));
  AND      g1486(.a(new_n999_), .b(i_2_5_148_0), .O(new_n1503_));
  AND      g1487(.a(new_n1503_), .b(new_n161_), .O(new_n1504_));
  AND      g1488(.a(new_n1382_), .b(new_n1158_), .O(new_n1505_));
  AND      g1489(.a(new_n1505_), .b(new_n1252_), .O(new_n1506_));
  OR       g1490(.a(new_n1506_), .b(new_n1504_), .O(new_n1507_));
  AND      g1491(.a(new_n1507_), .b(new_n20_), .O(new_n1508_));
  OR       g1492(.a(new_n1508_), .b(new_n1502_), .O(new_n1509_));
  OR       g1493(.a(new_n1509_), .b(new_n1479_), .O(new_n1510_));
  OR       g1494(.a(new_n1510_), .b(new_n1407_), .O(new_n1511_));
  AND      g1495(.a(new_n1511_), .b(i_2_5_102_0), .O(new_n1512_));
  OR       g1496(.a(i_2_5_84_0), .b(new_n221_), .O(new_n1513_));
  OR       g1497(.a(new_n1513_), .b(i_2_5_90_0), .O(new_n1514_));
  OR       g1498(.a(new_n1514_), .b(new_n27_), .O(new_n1515_));
  NAND     g1499(.a(new_n1515_), .b(new_n187_), .O(new_n1516_));
  AND      g1500(.a(new_n1516_), .b(new_n666_), .O(new_n1517_));
  OR       g1501(.a(new_n1517_), .b(new_n1041_), .O(new_n1518_));
  AND      g1502(.a(new_n1518_), .b(i_2_5_98_0), .O(new_n1519_));
  OR       g1503(.a(new_n1011_), .b(new_n319_), .O(new_n1520_));
  AND      g1504(.a(new_n1520_), .b(new_n21_), .O(new_n1521_));
  OR       g1505(.a(new_n1521_), .b(new_n79_), .O(new_n1522_));
  OR       g1506(.a(new_n1522_), .b(new_n1519_), .O(new_n1523_));
  AND      g1507(.a(new_n1523_), .b(i_2_5_62_0), .O(new_n1524_));
  AND      g1508(.a(new_n190_), .b(new_n21_), .O(new_n1525_));
  OR       g1509(.a(new_n1525_), .b(new_n1314_), .O(new_n1526_));
  OR       g1510(.a(new_n1526_), .b(new_n633_), .O(new_n1527_));
  AND      g1511(.a(new_n1527_), .b(i_2_5_62_0), .O(new_n1528_));
  NAND     g1512(.a(new_n40_), .b(new_n221_), .O(new_n1529_));
  AND      g1513(.a(new_n1529_), .b(i_2_5_148_0), .O(new_n1530_));
  AND      g1514(.a(new_n190_), .b(i_2_5_84_0), .O(new_n1531_));
  OR       g1515(.a(new_n1199_), .b(new_n326_), .O(new_n1532_));
  NAND     g1516(.a(new_n1532_), .b(new_n99_), .O(new_n1533_));
  AND      g1517(.a(new_n1533_), .b(new_n1531_), .O(new_n1534_));
  OR       g1518(.a(new_n1534_), .b(new_n1530_), .O(new_n1535_));
  OR       g1519(.a(new_n1535_), .b(new_n1528_), .O(new_n1536_));
  AND      g1520(.a(new_n1536_), .b(new_n19_), .O(new_n1537_));
  OR       g1521(.a(new_n822_), .b(i_2_5_90_0), .O(new_n1538_));
  OR       g1522(.a(new_n445_), .b(i_2_5_82_0), .O(new_n1539_));
  OR       g1523(.a(new_n1539_), .b(new_n1531_), .O(new_n1540_));
  NAND     g1524(.a(new_n279_), .b(i_2_5_98_0), .O(new_n1541_));
  AND      g1525(.a(new_n1541_), .b(new_n25_), .O(new_n1542_));
  NAND     g1526(.a(new_n1542_), .b(new_n1540_), .O(new_n1543_));
  NAND     g1527(.a(new_n1543_), .b(new_n1538_), .O(new_n1544_));
  OR       g1528(.a(new_n1544_), .b(new_n1537_), .O(new_n1545_));
  OR       g1529(.a(new_n1545_), .b(new_n1524_), .O(new_n1546_));
  AND      g1530(.a(new_n1546_), .b(new_n67_), .O(new_n1547_));
  AND      g1531(.a(i_2_5_82_0), .b(i_2_5_70_0), .O(new_n1548_));
  AND      g1532(.a(i_2_5_98_0), .b(i_2_5_70_0), .O(new_n1549_));
  AND      g1533(.a(new_n1549_), .b(new_n1394_), .O(new_n1550_));
  OR       g1534(.a(new_n1550_), .b(new_n1002_), .O(new_n1551_));
  AND      g1535(.a(new_n1551_), .b(i_2_5_42_0), .O(new_n1552_));
  OR       g1536(.a(new_n1552_), .b(new_n1548_), .O(new_n1553_));
  AND      g1537(.a(new_n1553_), .b(i_2_5_148_0), .O(new_n1554_));
  OR       g1538(.a(new_n261_), .b(new_n161_), .O(new_n1555_));
  AND      g1539(.a(new_n1555_), .b(new_n606_), .O(new_n1556_));
  AND      g1540(.a(new_n1059_), .b(new_n215_), .O(new_n1557_));
  OR       g1541(.a(new_n276_), .b(new_n28_), .O(new_n1558_));
  AND      g1542(.a(new_n1558_), .b(new_n99_), .O(new_n1559_));
  OR       g1543(.a(new_n1559_), .b(new_n1557_), .O(new_n1560_));
  OR       g1544(.a(new_n1560_), .b(new_n1556_), .O(new_n1561_));
  AND      g1545(.a(new_n1561_), .b(new_n21_), .O(new_n1562_));
  OR       g1546(.a(new_n261_), .b(new_n124_), .O(new_n1563_));
  AND      g1547(.a(new_n1563_), .b(i_2_5_12_0), .O(new_n1564_));
  OR       g1548(.a(new_n1564_), .b(new_n713_), .O(new_n1565_));
  OR       g1549(.a(new_n1565_), .b(new_n1562_), .O(new_n1566_));
  OR       g1550(.a(new_n1566_), .b(new_n1554_), .O(new_n1567_));
  AND      g1551(.a(new_n1567_), .b(new_n27_), .O(new_n1568_));
  AND      g1552(.a(new_n1054_), .b(new_n1002_), .O(new_n1569_));
  AND      g1553(.a(new_n1445_), .b(i_2_5_12_0), .O(new_n1570_));
  AND      g1554(.a(new_n261_), .b(new_n118_), .O(new_n1571_));
  OR       g1555(.a(new_n1571_), .b(new_n1570_), .O(new_n1572_));
  AND      g1556(.a(new_n1572_), .b(i_2_5_84_0), .O(new_n1573_));
  AND      g1557(.a(new_n319_), .b(new_n261_), .O(new_n1574_));
  OR       g1558(.a(new_n1574_), .b(new_n1573_), .O(new_n1575_));
  AND      g1559(.a(new_n1575_), .b(new_n21_), .O(new_n1576_));
  OR       g1560(.a(new_n1576_), .b(new_n1569_), .O(new_n1577_));
  OR       g1561(.a(new_n1577_), .b(new_n1568_), .O(new_n1578_));
  OR       g1562(.a(new_n1578_), .b(new_n1547_), .O(new_n1579_));
  AND      g1563(.a(new_n1579_), .b(new_n20_), .O(new_n1580_));
  OR       g1564(.a(new_n1360_), .b(new_n838_), .O(new_n1581_));
  AND      g1565(.a(new_n1581_), .b(i_2_5_12_0), .O(new_n1582_));
  OR       g1566(.a(new_n1372_), .b(new_n100_), .O(new_n1583_));
  AND      g1567(.a(new_n1583_), .b(new_n947_), .O(new_n1584_));
  OR       g1568(.a(new_n1584_), .b(new_n1582_), .O(new_n1585_));
  AND      g1569(.a(new_n1585_), .b(i_2_5_84_0), .O(new_n1586_));
  AND      g1570(.a(new_n838_), .b(new_n149_), .O(new_n1587_));
  OR       g1571(.a(new_n1587_), .b(new_n1586_), .O(new_n1588_));
  NAND     g1572(.a(new_n1588_), .b(new_n67_), .O(new_n1589_));
  NAND     g1573(.a(new_n33_), .b(i_2_5_12_0), .O(new_n1590_));
  OR       g1574(.a(new_n1590_), .b(new_n199_), .O(new_n1591_));
  NAND     g1575(.a(new_n1591_), .b(new_n1589_), .O(new_n1592_));
  AND      g1576(.a(new_n1592_), .b(new_n27_), .O(new_n1593_));
  OR       g1577(.a(new_n1392_), .b(new_n644_), .O(new_n1594_));
  NOT      g1578(.a(new_n1594_), .O(new_n1595_));
  AND      g1579(.a(new_n1595_), .b(new_n1002_), .O(new_n1596_));
  NOT      g1580(.a(new_n1161_), .O(new_n1597_));
  AND      g1581(.a(new_n1597_), .b(new_n45_), .O(new_n1598_));
  NOT      g1582(.a(new_n178_), .O(new_n1599_));
  NAND     g1583(.a(new_n1599_), .b(new_n68_), .O(new_n1600_));
  AND      g1584(.a(new_n1383_), .b(i_2_5_12_0), .O(new_n1601_));
  AND      g1585(.a(new_n1601_), .b(new_n1600_), .O(new_n1602_));
  OR       g1586(.a(new_n1602_), .b(new_n1598_), .O(new_n1603_));
  AND      g1587(.a(new_n1603_), .b(new_n19_), .O(new_n1604_));
  OR       g1588(.a(new_n1397_), .b(new_n199_), .O(new_n1605_));
  NAND     g1589(.a(new_n1605_), .b(i_2_5_70_0), .O(new_n1606_));
  NAND     g1590(.a(new_n1161_), .b(new_n112_), .O(new_n1607_));
  AND      g1591(.a(new_n1607_), .b(new_n45_), .O(new_n1608_));
  AND      g1592(.a(new_n1608_), .b(new_n1606_), .O(new_n1609_));
  OR       g1593(.a(new_n1609_), .b(new_n1604_), .O(new_n1610_));
  AND      g1594(.a(new_n1610_), .b(i_2_5_82_0), .O(new_n1611_));
  AND      g1595(.a(new_n1395_), .b(new_n838_), .O(new_n1612_));
  NOT      g1596(.a(new_n686_), .O(new_n1613_));
  AND      g1597(.a(new_n1598_), .b(new_n1613_), .O(new_n1614_));
  NOT      g1598(.a(new_n1360_), .O(new_n1615_));
  NAND     g1599(.a(new_n1454_), .b(new_n1615_), .O(new_n1616_));
  AND      g1600(.a(new_n1616_), .b(new_n645_), .O(new_n1617_));
  OR       g1601(.a(new_n1617_), .b(new_n1614_), .O(new_n1618_));
  AND      g1602(.a(new_n1618_), .b(i_2_5_84_0), .O(new_n1619_));
  OR       g1603(.a(new_n1619_), .b(new_n1612_), .O(new_n1620_));
  OR       g1604(.a(new_n1620_), .b(new_n1611_), .O(new_n1621_));
  AND      g1605(.a(new_n1621_), .b(i_2_5_42_0), .O(new_n1622_));
  OR       g1606(.a(new_n1622_), .b(new_n1596_), .O(new_n1623_));
  OR       g1607(.a(new_n1623_), .b(new_n1593_), .O(new_n1624_));
  OR       g1608(.a(new_n1624_), .b(new_n1580_), .O(new_n1625_));
  OR       g1609(.a(new_n1625_), .b(new_n1512_), .O(new_n1626_));
  AND      g1610(.a(new_n1626_), .b(new_n18_), .O(new_n1627_));
  NAND     g1611(.a(i_2_5_93_0), .b(i_2_5_90_0), .O(new_n1628_));
  OR       g1612(.a(new_n1628_), .b(new_n143_), .O(new_n1629_));
  OR       g1613(.a(i_2_5_90_0), .b(new_n99_), .O(new_n1630_));
  AND      g1614(.a(new_n1630_), .b(new_n130_), .O(new_n1631_));
  OR       g1615(.a(new_n1631_), .b(new_n221_), .O(new_n1632_));
  NAND     g1616(.a(new_n1632_), .b(new_n1629_), .O(new_n1633_));
  AND      g1617(.a(new_n1633_), .b(new_n51_), .O(new_n1634_));
  AND      g1618(.a(new_n118_), .b(new_n41_), .O(new_n1635_));
  AND      g1619(.a(new_n1419_), .b(new_n34_), .O(new_n1636_));
  OR       g1620(.a(new_n33_), .b(i_2_5_42_0), .O(new_n1637_));
  OR       g1621(.a(new_n1637_), .b(new_n1636_), .O(new_n1638_));
  AND      g1622(.a(new_n1638_), .b(i_2_5_62_0), .O(new_n1639_));
  OR       g1623(.a(new_n1639_), .b(new_n1635_), .O(new_n1640_));
  AND      g1624(.a(new_n1640_), .b(i_2_5_12_0), .O(new_n1641_));
  AND      g1625(.a(new_n1314_), .b(new_n198_), .O(new_n1642_));
  AND      g1626(.a(new_n244_), .b(new_n23_), .O(new_n1643_));
  NOT      g1627(.a(new_n31_), .O(new_n1644_));
  AND      g1628(.a(new_n319_), .b(new_n1644_), .O(new_n1645_));
  OR       g1629(.a(new_n1645_), .b(new_n1643_), .O(new_n1646_));
  AND      g1630(.a(new_n1646_), .b(new_n27_), .O(new_n1647_));
  OR       g1631(.a(new_n1647_), .b(new_n1642_), .O(new_n1648_));
  OR       g1632(.a(new_n1648_), .b(new_n1641_), .O(new_n1649_));
  AND      g1633(.a(new_n1649_), .b(new_n20_), .O(new_n1650_));
  OR       g1634(.a(new_n1650_), .b(new_n1634_), .O(new_n1651_));
  AND      g1635(.a(new_n1651_), .b(new_n19_), .O(new_n1652_));
  AND      g1636(.a(new_n456_), .b(new_n112_), .O(new_n1653_));
  OR       g1637(.a(new_n1653_), .b(new_n942_), .O(new_n1654_));
  NAND     g1638(.a(new_n1654_), .b(new_n797_), .O(new_n1655_));
  AND      g1639(.a(new_n1655_), .b(new_n27_), .O(new_n1656_));
  OR       g1640(.a(new_n998_), .b(i_2_5_99_0), .O(new_n1657_));
  OR       g1641(.a(new_n1657_), .b(new_n112_), .O(new_n1658_));
  NOT      g1642(.a(new_n1658_), .O(new_n1659_));
  OR       g1643(.a(new_n1659_), .b(new_n1656_), .O(new_n1660_));
  AND      g1644(.a(new_n1660_), .b(i_2_5_42_0), .O(new_n1661_));
  AND      g1645(.a(new_n998_), .b(i_2_5_99_0), .O(new_n1662_));
  NAND     g1646(.a(new_n1662_), .b(new_n1094_), .O(new_n1663_));
  AND      g1647(.a(new_n1663_), .b(new_n1058_), .O(new_n1664_));
  OR       g1648(.a(new_n1381_), .b(new_n20_), .O(new_n1665_));
  NAND     g1649(.a(new_n1630_), .b(new_n845_), .O(new_n1666_));
  AND      g1650(.a(new_n1666_), .b(new_n1665_), .O(new_n1667_));
  AND      g1651(.a(new_n1630_), .b(new_n810_), .O(new_n1668_));
  OR       g1652(.a(new_n1668_), .b(new_n130_), .O(new_n1669_));
  NAND     g1653(.a(new_n1669_), .b(new_n1657_), .O(new_n1670_));
  OR       g1654(.a(new_n1670_), .b(new_n1667_), .O(new_n1671_));
  OR       g1655(.a(new_n1671_), .b(new_n1664_), .O(new_n1672_));
  AND      g1656(.a(new_n1672_), .b(i_2_5_62_0), .O(new_n1673_));
  AND      g1657(.a(new_n1002_), .b(new_n278_), .O(new_n1674_));
  OR       g1658(.a(i_2_5_99_0), .b(new_n21_), .O(new_n1675_));
  OR       g1659(.a(new_n1675_), .b(new_n1493_), .O(new_n1676_));
  NAND     g1660(.a(new_n444_), .b(new_n45_), .O(new_n1677_));
  NAND     g1661(.a(new_n1677_), .b(new_n1676_), .O(new_n1678_));
  AND      g1662(.a(new_n1678_), .b(new_n99_), .O(new_n1679_));
  OR       g1663(.a(new_n1679_), .b(new_n1674_), .O(new_n1680_));
  OR       g1664(.a(new_n1680_), .b(new_n1673_), .O(new_n1681_));
  OR       g1665(.a(new_n1681_), .b(new_n1661_), .O(new_n1682_));
  AND      g1666(.a(new_n1682_), .b(i_2_5_148_0), .O(new_n1683_));
  OR       g1667(.a(new_n307_), .b(new_n732_), .O(new_n1684_));
  AND      g1668(.a(new_n1080_), .b(new_n20_), .O(new_n1685_));
  AND      g1669(.a(new_n1685_), .b(new_n1684_), .O(new_n1686_));
  NOT      g1670(.a(new_n871_), .O(new_n1687_));
  AND      g1671(.a(new_n380_), .b(i_2_5_12_0), .O(new_n1688_));
  AND      g1672(.a(new_n1688_), .b(new_n1687_), .O(new_n1689_));
  OR       g1673(.a(new_n1689_), .b(new_n1686_), .O(new_n1690_));
  AND      g1674(.a(new_n1690_), .b(new_n21_), .O(new_n1691_));
  OR       g1675(.a(new_n1691_), .b(new_n1683_), .O(new_n1692_));
  OR       g1676(.a(new_n1692_), .b(new_n1652_), .O(new_n1693_));
  AND      g1677(.a(new_n1693_), .b(i_2_5_102_0), .O(new_n1694_));
  AND      g1678(.a(new_n458_), .b(i_2_5_90_0), .O(new_n1695_));
  OR       g1679(.a(new_n1695_), .b(new_n35_), .O(new_n1696_));
  AND      g1680(.a(new_n1696_), .b(new_n20_), .O(new_n1697_));
  AND      g1681(.a(new_n1085_), .b(new_n112_), .O(new_n1698_));
  OR       g1682(.a(new_n1698_), .b(new_n79_), .O(new_n1699_));
  AND      g1683(.a(new_n1699_), .b(new_n20_), .O(new_n1700_));
  OR       g1684(.a(new_n1628_), .b(new_n113_), .O(new_n1701_));
  NAND     g1685(.a(new_n1701_), .b(new_n154_), .O(new_n1702_));
  AND      g1686(.a(new_n1702_), .b(i_2_5_42_0), .O(new_n1703_));
  OR       g1687(.a(i_2_5_102_0), .b(new_n99_), .O(new_n1704_));
  OR       g1688(.a(new_n18_), .b(i_2_5_84_0), .O(new_n1705_));
  OR       g1689(.a(new_n1705_), .b(new_n1704_), .O(new_n1706_));
  NAND     g1690(.a(new_n1706_), .b(new_n154_), .O(new_n1707_));
  AND      g1691(.a(new_n1707_), .b(i_2_5_12_0), .O(new_n1708_));
  OR       g1692(.a(new_n1708_), .b(new_n1703_), .O(new_n1709_));
  OR       g1693(.a(new_n1709_), .b(new_n1700_), .O(new_n1710_));
  AND      g1694(.a(new_n1710_), .b(new_n19_), .O(new_n1711_));
  OR       g1695(.a(new_n1711_), .b(new_n1697_), .O(new_n1712_));
  AND      g1696(.a(new_n1712_), .b(i_2_5_148_0), .O(new_n1713_));
  NOT      g1697(.a(new_n1514_), .O(new_n1714_));
  AND      g1698(.a(new_n1714_), .b(new_n1386_), .O(new_n1715_));
  AND      g1699(.a(new_n967_), .b(new_n19_), .O(new_n1716_));
  AND      g1700(.a(new_n1716_), .b(new_n1296_), .O(new_n1717_));
  AND      g1701(.a(new_n1057_), .b(new_n397_), .O(new_n1718_));
  OR       g1702(.a(new_n1718_), .b(new_n1495_), .O(new_n1719_));
  OR       g1703(.a(new_n1719_), .b(new_n1717_), .O(new_n1720_));
  AND      g1704(.a(new_n1720_), .b(i_2_5_84_0), .O(new_n1721_));
  OR       g1705(.a(new_n1721_), .b(new_n1715_), .O(new_n1722_));
  AND      g1706(.a(new_n1722_), .b(new_n27_), .O(new_n1723_));
  OR       g1707(.a(new_n1723_), .b(new_n1713_), .O(new_n1724_));
  AND      g1708(.a(new_n1724_), .b(i_2_5_62_0), .O(new_n1725_));
  AND      g1709(.a(new_n1675_), .b(i_2_5_42_0), .O(new_n1726_));
  OR       g1710(.a(new_n1726_), .b(new_n499_), .O(new_n1727_));
  AND      g1711(.a(new_n1727_), .b(new_n785_), .O(new_n1728_));
  NOT      g1712(.a(new_n1151_), .O(new_n1729_));
  AND      g1713(.a(new_n1729_), .b(new_n1141_), .O(new_n1730_));
  OR       g1714(.a(new_n1730_), .b(new_n1728_), .O(new_n1731_));
  AND      g1715(.a(new_n1731_), .b(new_n444_), .O(new_n1732_));
  AND      g1716(.a(new_n852_), .b(new_n741_), .O(new_n1733_));
  AND      g1717(.a(new_n1733_), .b(new_n1503_), .O(new_n1734_));
  OR       g1718(.a(new_n1734_), .b(new_n1732_), .O(new_n1735_));
  OR       g1719(.a(new_n1735_), .b(new_n1725_), .O(new_n1736_));
  OR       g1720(.a(new_n1736_), .b(new_n1694_), .O(new_n1737_));
  AND      g1721(.a(new_n1737_), .b(new_n67_), .O(new_n1738_));
  NOT      g1722(.a(new_n1043_), .O(new_n1739_));
  OR       g1723(.a(new_n20_), .b(i_2_5_84_0), .O(new_n1740_));
  OR       g1724(.a(new_n1740_), .b(new_n1161_), .O(new_n1741_));
  NAND     g1725(.a(new_n1741_), .b(new_n520_), .O(new_n1742_));
  AND      g1726(.a(new_n1742_), .b(new_n380_), .O(new_n1743_));
  AND      g1727(.a(new_n947_), .b(new_n470_), .O(new_n1744_));
  OR       g1728(.a(new_n1744_), .b(new_n1743_), .O(new_n1745_));
  AND      g1729(.a(new_n1745_), .b(new_n1739_), .O(new_n1746_));
  NOT      g1730(.a(new_n222_), .O(new_n1747_));
  NAND     g1731(.a(new_n637_), .b(new_n534_), .O(new_n1748_));
  NAND     g1732(.a(new_n1748_), .b(new_n844_), .O(new_n1749_));
  AND      g1733(.a(new_n1749_), .b(new_n19_), .O(new_n1750_));
  AND      g1734(.a(new_n1191_), .b(new_n99_), .O(new_n1751_));
  OR       g1735(.a(new_n1751_), .b(new_n1750_), .O(new_n1752_));
  AND      g1736(.a(new_n1752_), .b(new_n1747_), .O(new_n1753_));
  AND      g1737(.a(new_n1351_), .b(new_n65_), .O(new_n1754_));
  AND      g1738(.a(new_n1754_), .b(new_n351_), .O(new_n1755_));
  OR       g1739(.a(new_n1755_), .b(new_n1753_), .O(new_n1756_));
  AND      g1740(.a(new_n1756_), .b(new_n21_), .O(new_n1757_));
  OR       g1741(.a(new_n1382_), .b(new_n51_), .O(new_n1758_));
  AND      g1742(.a(new_n1758_), .b(new_n466_), .O(new_n1759_));
  OR       g1743(.a(new_n815_), .b(i_2_5_82_0), .O(new_n1760_));
  NAND     g1744(.a(new_n1760_), .b(new_n113_), .O(new_n1761_));
  AND      g1745(.a(new_n1761_), .b(i_2_5_42_0), .O(new_n1762_));
  OR       g1746(.a(new_n902_), .b(new_n72_), .O(new_n1763_));
  OR       g1747(.a(new_n68_), .b(i_2_5_98_0), .O(new_n1764_));
  NAND     g1748(.a(new_n1764_), .b(new_n1763_), .O(new_n1765_));
  AND      g1749(.a(new_n1765_), .b(new_n99_), .O(new_n1766_));
  OR       g1750(.a(new_n1766_), .b(new_n1762_), .O(new_n1767_));
  OR       g1751(.a(new_n1767_), .b(new_n1759_), .O(new_n1768_));
  AND      g1752(.a(new_n1768_), .b(i_2_5_148_0), .O(new_n1769_));
  OR       g1753(.a(new_n1043_), .b(new_n170_), .O(new_n1770_));
  NAND     g1754(.a(new_n1234_), .b(i_2_5_12_0), .O(new_n1771_));
  AND      g1755(.a(new_n815_), .b(i_2_5_84_0), .O(new_n1772_));
  AND      g1756(.a(new_n113_), .b(new_n221_), .O(new_n1773_));
  OR       g1757(.a(new_n1773_), .b(new_n1772_), .O(new_n1774_));
  OR       g1758(.a(new_n1774_), .b(new_n1771_), .O(new_n1775_));
  NAND     g1759(.a(new_n1775_), .b(new_n1770_), .O(new_n1776_));
  OR       g1760(.a(new_n1776_), .b(new_n1769_), .O(new_n1777_));
  AND      g1761(.a(new_n1777_), .b(new_n21_), .O(new_n1778_));
  AND      g1762(.a(new_n351_), .b(new_n50_), .O(new_n1779_));
  OR       g1763(.a(new_n784_), .b(new_n21_), .O(new_n1780_));
  AND      g1764(.a(new_n1780_), .b(new_n187_), .O(new_n1781_));
  OR       g1765(.a(new_n1781_), .b(new_n130_), .O(new_n1782_));
  OR       g1766(.a(new_n822_), .b(i_2_5_98_0), .O(new_n1783_));
  NAND     g1767(.a(new_n1783_), .b(new_n1782_), .O(new_n1784_));
  AND      g1768(.a(new_n1784_), .b(new_n426_), .O(new_n1785_));
  OR       g1769(.a(new_n1785_), .b(new_n1779_), .O(new_n1786_));
  OR       g1770(.a(new_n1786_), .b(new_n1778_), .O(new_n1787_));
  AND      g1771(.a(new_n1787_), .b(i_2_5_62_0), .O(new_n1788_));
  OR       g1772(.a(new_n1788_), .b(new_n1757_), .O(new_n1789_));
  AND      g1773(.a(new_n1789_), .b(new_n20_), .O(new_n1790_));
  OR       g1774(.a(new_n1790_), .b(new_n1746_), .O(new_n1791_));
  OR       g1775(.a(new_n1791_), .b(new_n1738_), .O(new_n1792_));
  OR       g1776(.a(new_n1792_), .b(new_n1627_), .O(new_n1793_));
  AND      g1777(.a(new_n1793_), .b(new_n54_), .O(new_n1794_));
  AND      g1778(.a(new_n45_), .b(new_n20_), .O(new_n1795_));
  AND      g1779(.a(new_n1705_), .b(i_2_5_12_0), .O(new_n1796_));
  AND      g1780(.a(new_n18_), .b(i_2_5_84_0), .O(new_n1797_));
  OR       g1781(.a(new_n1797_), .b(new_n319_), .O(new_n1798_));
  AND      g1782(.a(new_n1798_), .b(new_n1796_), .O(new_n1799_));
  AND      g1783(.a(new_n713_), .b(new_n18_), .O(new_n1800_));
  OR       g1784(.a(new_n1800_), .b(new_n1799_), .O(new_n1801_));
  AND      g1785(.a(new_n1801_), .b(new_n1795_), .O(new_n1802_));
  NAND     g1786(.a(new_n178_), .b(new_n20_), .O(new_n1803_));
  OR       g1787(.a(i_2_5_93_0), .b(new_n17_), .O(new_n1804_));
  OR       g1788(.a(new_n1804_), .b(new_n1513_), .O(new_n1805_));
  NAND     g1789(.a(new_n1805_), .b(new_n1803_), .O(new_n1806_));
  AND      g1790(.a(new_n1806_), .b(i_2_5_12_0), .O(new_n1807_));
  OR       g1791(.a(new_n112_), .b(i_2_5_82_0), .O(new_n1808_));
  AND      g1792(.a(new_n1795_), .b(new_n1808_), .O(new_n1809_));
  OR       g1793(.a(new_n1809_), .b(new_n1807_), .O(new_n1810_));
  AND      g1794(.a(new_n1810_), .b(i_2_5_42_0), .O(new_n1811_));
  AND      g1795(.a(new_n18_), .b(i_2_5_12_0), .O(new_n1812_));
  AND      g1796(.a(new_n18_), .b(i_2_5_62_0), .O(new_n1813_));
  AND      g1797(.a(new_n1813_), .b(new_n887_), .O(new_n1814_));
  OR       g1798(.a(new_n1814_), .b(new_n1812_), .O(new_n1815_));
  AND      g1799(.a(new_n1815_), .b(new_n864_), .O(new_n1816_));
  OR       g1800(.a(new_n1813_), .b(new_n444_), .O(new_n1817_));
  AND      g1801(.a(new_n1817_), .b(new_n20_), .O(new_n1818_));
  AND      g1802(.a(new_n1812_), .b(new_n178_), .O(new_n1819_));
  OR       g1803(.a(new_n1819_), .b(new_n1818_), .O(new_n1820_));
  AND      g1804(.a(new_n1820_), .b(new_n78_), .O(new_n1821_));
  OR       g1805(.a(new_n1821_), .b(new_n1816_), .O(new_n1822_));
  OR       g1806(.a(new_n1822_), .b(new_n1811_), .O(new_n1823_));
  AND      g1807(.a(new_n1823_), .b(new_n21_), .O(new_n1824_));
  OR       g1808(.a(new_n1824_), .b(new_n1802_), .O(new_n1825_));
  AND      g1809(.a(new_n1825_), .b(new_n67_), .O(new_n1826_));
  AND      g1810(.a(new_n1286_), .b(i_2_5_84_0), .O(new_n1827_));
  OR       g1811(.a(new_n1827_), .b(new_n1796_), .O(new_n1828_));
  AND      g1812(.a(new_n1828_), .b(new_n380_), .O(new_n1829_));
  OR       g1813(.a(new_n31_), .b(i_2_5_62_0), .O(new_n1830_));
  OR       g1814(.a(i_2_5_93_0), .b(i_2_5_70_0), .O(new_n1831_));
  NOT      g1815(.a(new_n1831_), .O(new_n1832_));
  AND      g1816(.a(new_n1832_), .b(new_n1830_), .O(new_n1833_));
  OR       g1817(.a(new_n1833_), .b(new_n1829_), .O(new_n1834_));
  AND      g1818(.a(new_n1834_), .b(i_2_5_82_0), .O(new_n1835_));
  AND      g1819(.a(new_n1286_), .b(new_n444_), .O(new_n1836_));
  OR       g1820(.a(new_n1836_), .b(new_n1835_), .O(new_n1837_));
  AND      g1821(.a(new_n1837_), .b(new_n20_), .O(new_n1838_));
  AND      g1822(.a(new_n1819_), .b(new_n527_), .O(new_n1839_));
  OR       g1823(.a(new_n526_), .b(i_2_5_93_0), .O(new_n1840_));
  NAND     g1824(.a(new_n1840_), .b(new_n740_), .O(new_n1841_));
  AND      g1825(.a(new_n1841_), .b(i_2_5_62_0), .O(new_n1842_));
  AND      g1826(.a(new_n736_), .b(i_2_5_82_0), .O(new_n1843_));
  AND      g1827(.a(new_n1812_), .b(i_2_5_70_0), .O(new_n1844_));
  OR       g1828(.a(new_n1844_), .b(new_n1843_), .O(new_n1845_));
  OR       g1829(.a(new_n1845_), .b(new_n1842_), .O(new_n1846_));
  AND      g1830(.a(new_n1846_), .b(i_2_5_84_0), .O(new_n1847_));
  NAND     g1831(.a(new_n1347_), .b(new_n1335_), .O(new_n1848_));
  OR       g1832(.a(new_n1424_), .b(new_n740_), .O(new_n1849_));
  NAND     g1833(.a(new_n1849_), .b(new_n1848_), .O(new_n1850_));
  AND      g1834(.a(new_n1850_), .b(new_n1644_), .O(new_n1851_));
  AND      g1835(.a(new_n210_), .b(new_n18_), .O(new_n1852_));
  OR       g1836(.a(new_n1852_), .b(new_n1851_), .O(new_n1853_));
  OR       g1837(.a(new_n1853_), .b(new_n1847_), .O(new_n1854_));
  AND      g1838(.a(new_n1854_), .b(new_n21_), .O(new_n1855_));
  OR       g1839(.a(new_n1855_), .b(new_n1839_), .O(new_n1856_));
  OR       g1840(.a(new_n1856_), .b(new_n1838_), .O(new_n1857_));
  AND      g1841(.a(new_n1857_), .b(new_n27_), .O(new_n1858_));
  AND      g1842(.a(new_n891_), .b(new_n221_), .O(new_n1859_));
  OR       g1843(.a(new_n1859_), .b(new_n432_), .O(new_n1860_));
  AND      g1844(.a(new_n1860_), .b(new_n20_), .O(new_n1861_));
  NAND     g1845(.a(new_n1514_), .b(new_n1808_), .O(new_n1862_));
  AND      g1846(.a(new_n1862_), .b(i_2_5_42_0), .O(new_n1863_));
  OR       g1847(.a(new_n1863_), .b(new_n1861_), .O(new_n1864_));
  AND      g1848(.a(new_n1864_), .b(new_n18_), .O(new_n1865_));
  AND      g1849(.a(new_n1063_), .b(i_2_5_12_0), .O(new_n1866_));
  OR       g1850(.a(i_2_5_93_0), .b(i_2_5_82_0), .O(new_n1867_));
  OR       g1851(.a(new_n1705_), .b(new_n130_), .O(new_n1868_));
  NAND     g1852(.a(new_n1868_), .b(new_n1867_), .O(new_n1869_));
  AND      g1853(.a(new_n1869_), .b(i_2_5_65_0), .O(new_n1870_));
  OR       g1854(.a(new_n1870_), .b(new_n1866_), .O(new_n1871_));
  AND      g1855(.a(new_n1871_), .b(new_n20_), .O(new_n1872_));
  OR       g1856(.a(new_n1872_), .b(new_n1865_), .O(new_n1873_));
  AND      g1857(.a(new_n1873_), .b(i_2_5_62_0), .O(new_n1874_));
  NAND     g1858(.a(new_n646_), .b(i_2_5_93_0), .O(new_n1875_));
  OR       g1859(.a(new_n1085_), .b(new_n20_), .O(new_n1876_));
  AND      g1860(.a(new_n1876_), .b(new_n444_), .O(new_n1877_));
  AND      g1861(.a(new_n1877_), .b(new_n1875_), .O(new_n1878_));
  OR       g1862(.a(new_n1878_), .b(new_n1874_), .O(new_n1879_));
  AND      g1863(.a(new_n1879_), .b(new_n67_), .O(new_n1880_));
  NAND     g1864(.a(new_n118_), .b(new_n112_), .O(new_n1881_));
  AND      g1865(.a(new_n500_), .b(i_2_5_12_0), .O(new_n1882_));
  OR       g1866(.a(i_2_5_99_0), .b(i_2_5_93_0), .O(new_n1883_));
  NOT      g1867(.a(new_n1883_), .O(new_n1884_));
  AND      g1868(.a(new_n1884_), .b(new_n1882_), .O(new_n1885_));
  AND      g1869(.a(new_n1885_), .b(new_n1881_), .O(new_n1886_));
  OR       g1870(.a(new_n1886_), .b(new_n1880_), .O(new_n1887_));
  OR       g1871(.a(new_n1887_), .b(new_n1858_), .O(new_n1888_));
  AND      g1872(.a(new_n1888_), .b(i_2_5_148_0), .O(new_n1889_));
  OR       g1873(.a(new_n1889_), .b(new_n1826_), .O(new_n1890_));
  AND      g1874(.a(new_n1890_), .b(new_n19_), .O(new_n1891_));
  AND      g1875(.a(new_n24_), .b(i_2_5_148_0), .O(new_n1892_));
  OR       g1876(.a(new_n1892_), .b(i_2_5_12_0), .O(new_n1893_));
  AND      g1877(.a(new_n1251_), .b(new_n67_), .O(new_n1894_));
  AND      g1878(.a(new_n1894_), .b(new_n1893_), .O(new_n1895_));
  AND      g1879(.a(new_n21_), .b(i_2_5_42_0), .O(new_n1896_));
  AND      g1880(.a(new_n1896_), .b(new_n1548_), .O(new_n1897_));
  OR       g1881(.a(new_n1882_), .b(new_n1046_), .O(new_n1898_));
  AND      g1882(.a(new_n1898_), .b(i_2_5_84_0), .O(new_n1899_));
  OR       g1883(.a(new_n1899_), .b(new_n1897_), .O(new_n1900_));
  OR       g1884(.a(new_n1900_), .b(new_n1895_), .O(new_n1901_));
  AND      g1885(.a(new_n1901_), .b(new_n27_), .O(new_n1902_));
  AND      g1886(.a(new_n1393_), .b(new_n624_), .O(new_n1903_));
  OR       g1887(.a(new_n1903_), .b(new_n1902_), .O(new_n1904_));
  AND      g1888(.a(new_n1904_), .b(i_2_5_62_0), .O(new_n1905_));
  OR       g1889(.a(new_n33_), .b(new_n67_), .O(new_n1906_));
  AND      g1890(.a(new_n1906_), .b(new_n458_), .O(new_n1907_));
  AND      g1891(.a(new_n1525_), .b(new_n527_), .O(new_n1908_));
  OR       g1892(.a(new_n1908_), .b(new_n1907_), .O(new_n1909_));
  AND      g1893(.a(new_n1909_), .b(i_2_5_84_0), .O(new_n1910_));
  OR       g1894(.a(new_n1910_), .b(new_n1595_), .O(new_n1911_));
  OR       g1895(.a(new_n1911_), .b(new_n1905_), .O(new_n1912_));
  AND      g1896(.a(new_n1912_), .b(new_n18_), .O(new_n1913_));
  OR       g1897(.a(new_n1594_), .b(new_n221_), .O(new_n1914_));
  NOT      g1898(.a(new_n1424_), .O(new_n1915_));
  AND      g1899(.a(new_n22_), .b(i_2_5_148_0), .O(new_n1916_));
  AND      g1900(.a(new_n1916_), .b(new_n1915_), .O(new_n1917_));
  NAND     g1901(.a(new_n1590_), .b(new_n519_), .O(new_n1918_));
  AND      g1902(.a(new_n1918_), .b(new_n30_), .O(new_n1919_));
  OR       g1903(.a(new_n1919_), .b(new_n1917_), .O(new_n1920_));
  NAND     g1904(.a(new_n1920_), .b(new_n380_), .O(new_n1921_));
  NAND     g1905(.a(new_n1921_), .b(new_n1914_), .O(new_n1922_));
  OR       g1906(.a(new_n1922_), .b(new_n1913_), .O(new_n1923_));
  AND      g1907(.a(new_n1923_), .b(new_n20_), .O(new_n1924_));
  NAND     g1908(.a(new_n961_), .b(new_n444_), .O(new_n1925_));
  OR       g1909(.a(new_n1740_), .b(new_n474_), .O(new_n1926_));
  OR       g1910(.a(new_n1926_), .b(new_n1099_), .O(new_n1927_));
  NAND     g1911(.a(new_n1927_), .b(new_n1925_), .O(new_n1928_));
  AND      g1912(.a(new_n1393_), .b(new_n45_), .O(new_n1929_));
  AND      g1913(.a(new_n1929_), .b(new_n1928_), .O(new_n1930_));
  OR       g1914(.a(new_n1930_), .b(new_n1924_), .O(new_n1931_));
  OR       g1915(.a(new_n1931_), .b(new_n1891_), .O(new_n1932_));
  AND      g1916(.a(new_n1932_), .b(i_2_5_102_0), .O(new_n1933_));
  OR       g1917(.a(new_n1896_), .b(new_n444_), .O(new_n1934_));
  AND      g1918(.a(new_n1934_), .b(new_n785_), .O(new_n1935_));
  OR       g1919(.a(new_n1178_), .b(new_n19_), .O(new_n1936_));
  NAND     g1920(.a(new_n1936_), .b(new_n32_), .O(new_n1937_));
  NAND     g1921(.a(new_n1937_), .b(new_n1199_), .O(new_n1938_));
  AND      g1922(.a(new_n1938_), .b(i_2_5_82_0), .O(new_n1939_));
  OR       g1923(.a(new_n1939_), .b(new_n1935_), .O(new_n1940_));
  AND      g1924(.a(new_n1940_), .b(new_n67_), .O(new_n1941_));
  OR       g1925(.a(new_n713_), .b(new_n21_), .O(new_n1942_));
  AND      g1926(.a(new_n1942_), .b(new_n27_), .O(new_n1943_));
  NAND     g1927(.a(i_2_5_70_0), .b(i_2_5_65_0), .O(new_n1944_));
  OR       g1928(.a(new_n1944_), .b(new_n550_), .O(new_n1945_));
  NAND     g1929(.a(new_n1945_), .b(i_2_5_90_0), .O(new_n1946_));
  AND      g1930(.a(new_n1946_), .b(i_2_5_42_0), .O(new_n1947_));
  OR       g1931(.a(new_n1947_), .b(new_n1943_), .O(new_n1948_));
  AND      g1932(.a(new_n1948_), .b(i_2_5_12_0), .O(new_n1949_));
  AND      g1933(.a(new_n999_), .b(new_n713_), .O(new_n1950_));
  OR       g1934(.a(new_n1950_), .b(new_n1949_), .O(new_n1951_));
  OR       g1935(.a(new_n1951_), .b(new_n1941_), .O(new_n1952_));
  AND      g1936(.a(new_n1952_), .b(i_2_5_148_0), .O(new_n1953_));
  OR       g1937(.a(new_n444_), .b(new_n319_), .O(new_n1954_));
  OR       g1938(.a(new_n1392_), .b(new_n784_), .O(new_n1955_));
  NOT      g1939(.a(new_n1955_), .O(new_n1956_));
  AND      g1940(.a(new_n1956_), .b(new_n1954_), .O(new_n1957_));
  OR       g1941(.a(new_n1957_), .b(new_n1953_), .O(new_n1958_));
  AND      g1942(.a(new_n1958_), .b(new_n20_), .O(new_n1959_));
  NAND     g1943(.a(new_n552_), .b(i_2_5_90_0), .O(new_n1960_));
  NOT      g1944(.a(new_n1455_), .O(new_n1961_));
  AND      g1945(.a(new_n1961_), .b(new_n1351_), .O(new_n1962_));
  AND      g1946(.a(new_n1962_), .b(new_n1960_), .O(new_n1963_));
  OR       g1947(.a(new_n1963_), .b(new_n1959_), .O(new_n1964_));
  AND      g1948(.a(new_n1964_), .b(new_n18_), .O(new_n1965_));
  NOT      g1949(.a(new_n1028_), .O(new_n1966_));
  OR       g1950(.a(new_n1191_), .b(new_n1966_), .O(new_n1967_));
  AND      g1951(.a(new_n1967_), .b(new_n458_), .O(new_n1968_));
  NOT      g1952(.a(new_n1460_), .O(new_n1969_));
  AND      g1953(.a(new_n1916_), .b(new_n1969_), .O(new_n1970_));
  OR       g1954(.a(new_n1970_), .b(new_n1968_), .O(new_n1971_));
  OR       g1955(.a(new_n810_), .b(i_2_5_70_0), .O(new_n1972_));
  NOT      g1956(.a(new_n1972_), .O(new_n1973_));
  AND      g1957(.a(new_n1973_), .b(new_n1971_), .O(new_n1974_));
  OR       g1958(.a(new_n1974_), .b(new_n1965_), .O(new_n1975_));
  AND      g1959(.a(new_n1975_), .b(i_2_5_62_0), .O(new_n1976_));
  OR       g1960(.a(new_n735_), .b(new_n279_), .O(new_n1977_));
  NAND     g1961(.a(new_n1977_), .b(new_n1532_), .O(new_n1978_));
  AND      g1962(.a(new_n1978_), .b(new_n838_), .O(new_n1979_));
  NAND     g1963(.a(new_n1704_), .b(new_n747_), .O(new_n1980_));
  AND      g1964(.a(new_n1944_), .b(i_2_5_82_0), .O(new_n1981_));
  AND      g1965(.a(new_n1981_), .b(new_n196_), .O(new_n1982_));
  AND      g1966(.a(new_n1982_), .b(new_n1980_), .O(new_n1983_));
  OR       g1967(.a(new_n1983_), .b(new_n1979_), .O(new_n1984_));
  AND      g1968(.a(new_n1984_), .b(new_n1812_), .O(new_n1985_));
  OR       g1969(.a(new_n1985_), .b(new_n1976_), .O(new_n1986_));
  OR       g1970(.a(new_n1986_), .b(new_n1933_), .O(new_n1987_));
  OR       g1971(.a(new_n1987_), .b(new_n1794_), .O(new_n1988_));
  OR       g1972(.a(new_n1988_), .b(new_n1346_), .O(o_2_5_0_0));
endmodule


