// Benchmark "kernel_2_6" written by ABC on Wed May  4 18:34:14 2022

module kernel_2_6 ( 
    i_2_6_5_0, i_2_6_32_0, i_2_6_33_0, i_2_6_34_0, i_2_6_40_0, i_2_6_51_0,
    i_2_6_62_0, i_2_6_63_0, i_2_6_84_0, i_2_6_110_0, i_2_6_111_0,
    i_2_6_118_0, i_2_6_120_0, i_2_6_124_0, i_2_6_142_0,
    o_2_6_0_0  );
  input  i_2_6_5_0, i_2_6_32_0, i_2_6_33_0, i_2_6_34_0, i_2_6_40_0,
    i_2_6_51_0, i_2_6_62_0, i_2_6_63_0, i_2_6_84_0, i_2_6_110_0,
    i_2_6_111_0, i_2_6_118_0, i_2_6_120_0, i_2_6_124_0, i_2_6_142_0;
  output o_2_6_0_0;
  wire new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_;
  NOT      g0000(.a(i_2_6_120_0), .O(new_n17_));
  NOT      g0001(.a(i_2_6_118_0), .O(new_n18_));
  NOT      g0002(.a(i_2_6_124_0), .O(new_n19_));
  NOT      g0003(.a(i_2_6_110_0), .O(new_n20_));
  NOT      g0004(.a(i_2_6_32_0), .O(new_n21_));
  NOT      g0005(.a(i_2_6_111_0), .O(new_n22_));
  NOT      g0006(.a(i_2_6_40_0), .O(new_n23_));
  OR       g0007(.a(i_2_6_142_0), .b(new_n23_), .O(new_n24_));
  OR       g0008(.a(new_n24_), .b(new_n22_), .O(new_n25_));
  NOT      g0009(.a(i_2_6_62_0), .O(new_n26_));
  OR       g0010(.a(i_2_6_84_0), .b(new_n26_), .O(new_n27_));
  NOT      g0011(.a(i_2_6_142_0), .O(new_n28_));
  OR       g0012(.a(i_2_6_63_0), .b(i_2_6_40_0), .O(new_n29_));
  OR       g0013(.a(new_n29_), .b(new_n28_), .O(new_n30_));
  OR       g0014(.a(new_n30_), .b(new_n27_), .O(new_n31_));
  NAND     g0015(.a(new_n31_), .b(new_n25_), .O(new_n32_));
  AND      g0016(.a(new_n32_), .b(new_n21_), .O(new_n33_));
  AND      g0017(.a(i_2_6_111_0), .b(i_2_6_32_0), .O(new_n34_));
  NOT      g0018(.a(i_2_6_84_0), .O(new_n35_));
  AND      g0019(.a(new_n35_), .b(i_2_6_63_0), .O(new_n36_));
  AND      g0020(.a(new_n36_), .b(new_n34_), .O(new_n37_));
  OR       g0021(.a(new_n37_), .b(new_n33_), .O(new_n38_));
  AND      g0022(.a(new_n38_), .b(new_n20_), .O(new_n39_));
  AND      g0023(.a(i_2_6_34_0), .b(i_2_6_32_0), .O(new_n40_));
  AND      g0024(.a(new_n35_), .b(i_2_6_32_0), .O(new_n41_));
  OR       g0025(.a(new_n41_), .b(i_2_6_34_0), .O(new_n42_));
  AND      g0026(.a(new_n42_), .b(i_2_6_63_0), .O(new_n43_));
  OR       g0027(.a(new_n43_), .b(new_n40_), .O(new_n44_));
  AND      g0028(.a(new_n44_), .b(i_2_6_142_0), .O(new_n45_));
  AND      g0029(.a(i_2_6_110_0), .b(new_n35_), .O(new_n46_));
  OR       g0030(.a(new_n46_), .b(i_2_6_111_0), .O(new_n47_));
  NAND     g0031(.a(new_n47_), .b(i_2_6_34_0), .O(new_n48_));
  NAND     g0032(.a(i_2_6_51_0), .b(i_2_6_32_0), .O(new_n49_));
  OR       g0033(.a(i_2_6_142_0), .b(new_n20_), .O(new_n50_));
  OR       g0034(.a(new_n50_), .b(new_n22_), .O(new_n51_));
  OR       g0035(.a(new_n51_), .b(new_n49_), .O(new_n52_));
  NAND     g0036(.a(new_n52_), .b(new_n48_), .O(new_n53_));
  OR       g0037(.a(new_n53_), .b(new_n45_), .O(new_n54_));
  AND      g0038(.a(new_n54_), .b(new_n23_), .O(new_n55_));
  OR       g0039(.a(i_2_6_110_0), .b(i_2_6_63_0), .O(new_n56_));
  AND      g0040(.a(new_n56_), .b(new_n40_), .O(new_n57_));
  AND      g0041(.a(i_2_6_142_0), .b(i_2_6_111_0), .O(new_n58_));
  AND      g0042(.a(new_n58_), .b(i_2_6_63_0), .O(new_n59_));
  AND      g0043(.a(new_n59_), .b(i_2_6_51_0), .O(new_n60_));
  OR       g0044(.a(new_n60_), .b(new_n57_), .O(new_n61_));
  OR       g0045(.a(new_n61_), .b(new_n55_), .O(new_n62_));
  AND      g0046(.a(new_n62_), .b(i_2_6_62_0), .O(new_n63_));
  OR       g0047(.a(new_n63_), .b(new_n39_), .O(new_n64_));
  AND      g0048(.a(new_n64_), .b(new_n19_), .O(new_n65_));
  NAND     g0049(.a(i_2_6_110_0), .b(i_2_6_63_0), .O(new_n66_));
  NAND     g0050(.a(new_n66_), .b(i_2_6_40_0), .O(new_n67_));
  AND      g0051(.a(i_2_6_142_0), .b(i_2_6_110_0), .O(new_n68_));
  OR       g0052(.a(new_n68_), .b(i_2_6_63_0), .O(new_n69_));
  AND      g0053(.a(new_n69_), .b(i_2_6_62_0), .O(new_n70_));
  AND      g0054(.a(new_n70_), .b(new_n67_), .O(new_n71_));
  AND      g0055(.a(i_2_6_111_0), .b(i_2_6_63_0), .O(new_n72_));
  AND      g0056(.a(i_2_6_111_0), .b(new_n23_), .O(new_n73_));
  AND      g0057(.a(new_n73_), .b(i_2_6_110_0), .O(new_n74_));
  OR       g0058(.a(new_n74_), .b(new_n72_), .O(new_n75_));
  OR       g0059(.a(new_n75_), .b(new_n71_), .O(new_n76_));
  AND      g0060(.a(new_n76_), .b(i_2_6_32_0), .O(new_n77_));
  NOT      g0061(.a(new_n66_), .O(new_n78_));
  AND      g0062(.a(i_2_6_111_0), .b(new_n20_), .O(new_n79_));
  OR       g0063(.a(new_n79_), .b(new_n78_), .O(new_n80_));
  AND      g0064(.a(i_2_6_111_0), .b(i_2_6_110_0), .O(new_n81_));
  OR       g0065(.a(new_n81_), .b(new_n23_), .O(new_n82_));
  AND      g0066(.a(new_n82_), .b(i_2_6_62_0), .O(new_n83_));
  AND      g0067(.a(new_n83_), .b(new_n80_), .O(new_n84_));
  AND      g0068(.a(i_2_6_142_0), .b(i_2_6_32_0), .O(new_n85_));
  AND      g0069(.a(new_n85_), .b(new_n29_), .O(new_n86_));
  OR       g0070(.a(new_n86_), .b(new_n36_), .O(new_n87_));
  OR       g0071(.a(i_2_6_110_0), .b(new_n23_), .O(new_n88_));
  AND      g0072(.a(new_n88_), .b(new_n19_), .O(new_n89_));
  AND      g0073(.a(new_n89_), .b(new_n87_), .O(new_n90_));
  OR       g0074(.a(new_n90_), .b(new_n84_), .O(new_n91_));
  OR       g0075(.a(new_n91_), .b(new_n77_), .O(new_n92_));
  AND      g0076(.a(new_n92_), .b(i_2_6_34_0), .O(new_n93_));
  AND      g0077(.a(i_2_6_124_0), .b(i_2_6_40_0), .O(new_n94_));
  AND      g0078(.a(i_2_6_63_0), .b(new_n23_), .O(new_n95_));
  AND      g0079(.a(new_n95_), .b(i_2_6_62_0), .O(new_n96_));
  OR       g0080(.a(new_n96_), .b(new_n94_), .O(new_n97_));
  AND      g0081(.a(new_n97_), .b(i_2_6_32_0), .O(new_n98_));
  OR       g0082(.a(new_n95_), .b(i_2_6_142_0), .O(new_n99_));
  OR       g0083(.a(i_2_6_63_0), .b(i_2_6_62_0), .O(new_n100_));
  AND      g0084(.a(new_n100_), .b(i_2_6_34_0), .O(new_n101_));
  AND      g0085(.a(i_2_6_111_0), .b(i_2_6_62_0), .O(new_n102_));
  AND      g0086(.a(i_2_6_63_0), .b(i_2_6_40_0), .O(new_n103_));
  OR       g0087(.a(new_n103_), .b(new_n102_), .O(new_n104_));
  OR       g0088(.a(new_n104_), .b(new_n101_), .O(new_n105_));
  AND      g0089(.a(new_n105_), .b(new_n99_), .O(new_n106_));
  OR       g0090(.a(new_n106_), .b(new_n98_), .O(new_n107_));
  AND      g0091(.a(new_n107_), .b(i_2_6_110_0), .O(new_n108_));
  AND      g0092(.a(i_2_6_142_0), .b(new_n23_), .O(new_n109_));
  OR       g0093(.a(new_n109_), .b(i_2_6_62_0), .O(new_n110_));
  AND      g0094(.a(new_n110_), .b(i_2_6_63_0), .O(new_n111_));
  AND      g0095(.a(i_2_6_63_0), .b(i_2_6_32_0), .O(new_n112_));
  OR       g0096(.a(new_n112_), .b(i_2_6_111_0), .O(new_n113_));
  AND      g0097(.a(new_n23_), .b(i_2_6_32_0), .O(new_n114_));
  AND      g0098(.a(new_n114_), .b(i_2_6_62_0), .O(new_n115_));
  OR       g0099(.a(new_n115_), .b(new_n113_), .O(new_n116_));
  OR       g0100(.a(new_n116_), .b(new_n111_), .O(new_n117_));
  AND      g0101(.a(new_n117_), .b(i_2_6_34_0), .O(new_n118_));
  AND      g0102(.a(new_n114_), .b(new_n20_), .O(new_n119_));
  AND      g0103(.a(new_n119_), .b(new_n72_), .O(new_n120_));
  OR       g0104(.a(new_n120_), .b(new_n118_), .O(new_n121_));
  OR       g0105(.a(new_n121_), .b(new_n108_), .O(new_n122_));
  AND      g0106(.a(new_n122_), .b(new_n35_), .O(new_n123_));
  OR       g0107(.a(new_n123_), .b(new_n93_), .O(new_n124_));
  OR       g0108(.a(new_n124_), .b(new_n65_), .O(new_n125_));
  AND      g0109(.a(new_n125_), .b(new_n18_), .O(new_n126_));
  AND      g0110(.a(i_2_6_142_0), .b(new_n19_), .O(new_n127_));
  OR       g0111(.a(new_n127_), .b(new_n36_), .O(new_n128_));
  OR       g0112(.a(new_n35_), .b(i_2_6_63_0), .O(new_n129_));
  AND      g0113(.a(new_n129_), .b(new_n23_), .O(new_n130_));
  AND      g0114(.a(new_n130_), .b(new_n128_), .O(new_n131_));
  OR       g0115(.a(new_n95_), .b(new_n35_), .O(new_n132_));
  AND      g0116(.a(new_n132_), .b(i_2_6_111_0), .O(new_n133_));
  OR       g0117(.a(i_2_6_124_0), .b(i_2_6_84_0), .O(new_n134_));
  NOT      g0118(.a(new_n134_), .O(new_n135_));
  AND      g0119(.a(new_n135_), .b(i_2_6_63_0), .O(new_n136_));
  OR       g0120(.a(new_n136_), .b(new_n133_), .O(new_n137_));
  OR       g0121(.a(new_n137_), .b(new_n131_), .O(new_n138_));
  AND      g0122(.a(new_n138_), .b(i_2_6_32_0), .O(new_n139_));
  OR       g0123(.a(i_2_6_142_0), .b(new_n19_), .O(new_n140_));
  AND      g0124(.a(new_n140_), .b(new_n129_), .O(new_n141_));
  OR       g0125(.a(new_n141_), .b(new_n72_), .O(new_n142_));
  AND      g0126(.a(new_n142_), .b(i_2_6_32_0), .O(new_n143_));
  AND      g0127(.a(i_2_6_142_0), .b(i_2_6_63_0), .O(new_n144_));
  OR       g0128(.a(new_n144_), .b(new_n41_), .O(new_n145_));
  AND      g0129(.a(new_n145_), .b(i_2_6_40_0), .O(new_n146_));
  OR       g0130(.a(new_n146_), .b(new_n143_), .O(new_n147_));
  AND      g0131(.a(new_n147_), .b(i_2_6_110_0), .O(new_n148_));
  AND      g0132(.a(i_2_6_110_0), .b(new_n23_), .O(new_n149_));
  OR       g0133(.a(new_n127_), .b(i_2_6_111_0), .O(new_n150_));
  AND      g0134(.a(new_n150_), .b(new_n23_), .O(new_n151_));
  OR       g0135(.a(new_n151_), .b(new_n149_), .O(new_n152_));
  AND      g0136(.a(new_n152_), .b(new_n36_), .O(new_n153_));
  OR       g0137(.a(new_n153_), .b(new_n148_), .O(new_n154_));
  OR       g0138(.a(new_n154_), .b(new_n139_), .O(new_n155_));
  AND      g0139(.a(new_n155_), .b(i_2_6_62_0), .O(new_n156_));
  AND      g0140(.a(new_n140_), .b(i_2_6_110_0), .O(new_n157_));
  AND      g0141(.a(new_n73_), .b(new_n35_), .O(new_n158_));
  AND      g0142(.a(new_n158_), .b(new_n157_), .O(new_n159_));
  AND      g0143(.a(i_2_6_124_0), .b(new_n35_), .O(new_n160_));
  OR       g0144(.a(new_n160_), .b(i_2_6_142_0), .O(new_n161_));
  AND      g0145(.a(new_n161_), .b(new_n81_), .O(new_n162_));
  OR       g0146(.a(i_2_6_111_0), .b(new_n35_), .O(new_n163_));
  AND      g0147(.a(new_n163_), .b(i_2_6_142_0), .O(new_n164_));
  AND      g0148(.a(new_n164_), .b(new_n114_), .O(new_n165_));
  AND      g0149(.a(i_2_6_111_0), .b(new_n35_), .O(new_n166_));
  AND      g0150(.a(new_n166_), .b(i_2_6_32_0), .O(new_n167_));
  OR       g0151(.a(new_n73_), .b(new_n41_), .O(new_n168_));
  AND      g0152(.a(new_n168_), .b(i_2_6_110_0), .O(new_n169_));
  OR       g0153(.a(new_n169_), .b(new_n167_), .O(new_n170_));
  OR       g0154(.a(new_n170_), .b(new_n165_), .O(new_n171_));
  AND      g0155(.a(new_n171_), .b(new_n19_), .O(new_n172_));
  OR       g0156(.a(new_n172_), .b(new_n162_), .O(new_n173_));
  AND      g0157(.a(new_n173_), .b(i_2_6_63_0), .O(new_n174_));
  OR       g0158(.a(new_n174_), .b(new_n159_), .O(new_n175_));
  OR       g0159(.a(new_n175_), .b(new_n156_), .O(new_n176_));
  AND      g0160(.a(new_n176_), .b(i_2_6_34_0), .O(new_n177_));
  AND      g0161(.a(i_2_6_142_0), .b(new_n35_), .O(new_n178_));
  AND      g0162(.a(i_2_6_124_0), .b(i_2_6_110_0), .O(new_n179_));
  NOT      g0163(.a(new_n179_), .O(new_n180_));
  NAND     g0164(.a(new_n180_), .b(new_n178_), .O(new_n181_));
  AND      g0165(.a(i_2_6_142_0), .b(i_2_6_124_0), .O(new_n182_));
  NOT      g0166(.a(new_n182_), .O(new_n183_));
  AND      g0167(.a(new_n183_), .b(new_n134_), .O(new_n184_));
  NAND     g0168(.a(new_n114_), .b(i_2_6_110_0), .O(new_n185_));
  OR       g0169(.a(new_n185_), .b(new_n184_), .O(new_n186_));
  NAND     g0170(.a(new_n186_), .b(new_n181_), .O(new_n187_));
  AND      g0171(.a(new_n72_), .b(i_2_6_62_0), .O(new_n188_));
  AND      g0172(.a(new_n188_), .b(new_n187_), .O(new_n189_));
  OR       g0173(.a(new_n189_), .b(new_n177_), .O(new_n190_));
  OR       g0174(.a(new_n190_), .b(new_n126_), .O(new_n191_));
  AND      g0175(.a(new_n191_), .b(i_2_6_33_0), .O(new_n192_));
  NOT      g0176(.a(i_2_6_51_0), .O(new_n193_));
  AND      g0177(.a(new_n18_), .b(i_2_6_32_0), .O(new_n194_));
  AND      g0178(.a(i_2_6_110_0), .b(i_2_6_40_0), .O(new_n195_));
  AND      g0179(.a(new_n195_), .b(i_2_6_111_0), .O(new_n196_));
  OR       g0180(.a(new_n196_), .b(new_n194_), .O(new_n197_));
  AND      g0181(.a(new_n197_), .b(i_2_6_62_0), .O(new_n198_));
  AND      g0182(.a(new_n18_), .b(i_2_6_110_0), .O(new_n199_));
  AND      g0183(.a(new_n135_), .b(new_n79_), .O(new_n200_));
  OR       g0184(.a(new_n200_), .b(new_n199_), .O(new_n201_));
  AND      g0185(.a(new_n201_), .b(i_2_6_32_0), .O(new_n202_));
  OR       g0186(.a(new_n202_), .b(new_n198_), .O(new_n203_));
  AND      g0187(.a(new_n203_), .b(i_2_6_142_0), .O(new_n204_));
  OR       g0188(.a(i_2_6_118_0), .b(i_2_6_110_0), .O(new_n205_));
  NOT      g0189(.a(new_n205_), .O(new_n206_));
  OR       g0190(.a(new_n166_), .b(new_n34_), .O(new_n207_));
  AND      g0191(.a(new_n207_), .b(new_n206_), .O(new_n208_));
  OR       g0192(.a(new_n208_), .b(new_n204_), .O(new_n209_));
  AND      g0193(.a(new_n209_), .b(i_2_6_34_0), .O(new_n210_));
  AND      g0194(.a(i_2_6_142_0), .b(i_2_6_118_0), .O(new_n211_));
  AND      g0195(.a(new_n211_), .b(new_n19_), .O(new_n212_));
  OR       g0196(.a(new_n212_), .b(new_n41_), .O(new_n213_));
  NOT      g0197(.a(new_n94_), .O(new_n214_));
  AND      g0198(.a(new_n214_), .b(i_2_6_63_0), .O(new_n215_));
  AND      g0199(.a(new_n215_), .b(new_n213_), .O(new_n216_));
  AND      g0200(.a(new_n19_), .b(i_2_6_63_0), .O(new_n217_));
  AND      g0201(.a(new_n217_), .b(i_2_6_32_0), .O(new_n218_));
  OR       g0202(.a(new_n218_), .b(new_n160_), .O(new_n219_));
  AND      g0203(.a(new_n219_), .b(new_n18_), .O(new_n220_));
  AND      g0204(.a(i_2_6_124_0), .b(new_n20_), .O(new_n221_));
  OR       g0205(.a(new_n221_), .b(new_n35_), .O(new_n222_));
  NOT      g0206(.a(new_n160_), .O(new_n223_));
  AND      g0207(.a(new_n223_), .b(new_n109_), .O(new_n224_));
  AND      g0208(.a(new_n224_), .b(new_n222_), .O(new_n225_));
  OR       g0209(.a(new_n225_), .b(new_n220_), .O(new_n226_));
  OR       g0210(.a(new_n226_), .b(new_n216_), .O(new_n227_));
  AND      g0211(.a(new_n227_), .b(i_2_6_111_0), .O(new_n228_));
  OR       g0212(.a(i_2_6_124_0), .b(i_2_6_40_0), .O(new_n229_));
  NOT      g0213(.a(new_n229_), .O(new_n230_));
  AND      g0214(.a(new_n230_), .b(new_n163_), .O(new_n231_));
  OR       g0215(.a(new_n231_), .b(new_n167_), .O(new_n232_));
  AND      g0216(.a(new_n232_), .b(i_2_6_63_0), .O(new_n233_));
  OR       g0217(.a(i_2_6_111_0), .b(i_2_6_63_0), .O(new_n234_));
  NAND     g0218(.a(new_n234_), .b(new_n229_), .O(new_n235_));
  OR       g0219(.a(i_2_6_124_0), .b(i_2_6_63_0), .O(new_n236_));
  AND      g0220(.a(new_n236_), .b(i_2_6_32_0), .O(new_n237_));
  AND      g0221(.a(new_n237_), .b(new_n235_), .O(new_n238_));
  NOT      g0222(.a(i_2_6_63_0), .O(new_n239_));
  AND      g0223(.a(new_n182_), .b(new_n239_), .O(new_n240_));
  OR       g0224(.a(new_n240_), .b(new_n35_), .O(new_n241_));
  OR       g0225(.a(new_n241_), .b(new_n238_), .O(new_n242_));
  AND      g0226(.a(new_n242_), .b(new_n18_), .O(new_n243_));
  OR       g0227(.a(new_n243_), .b(new_n233_), .O(new_n244_));
  AND      g0228(.a(new_n244_), .b(i_2_6_110_0), .O(new_n245_));
  OR       g0229(.a(i_2_6_118_0), .b(i_2_6_40_0), .O(new_n246_));
  NOT      g0230(.a(new_n246_), .O(new_n247_));
  AND      g0231(.a(new_n247_), .b(i_2_6_142_0), .O(new_n248_));
  AND      g0232(.a(new_n248_), .b(new_n218_), .O(new_n249_));
  OR       g0233(.a(new_n249_), .b(new_n245_), .O(new_n250_));
  OR       g0234(.a(new_n250_), .b(new_n228_), .O(new_n251_));
  AND      g0235(.a(new_n251_), .b(i_2_6_62_0), .O(new_n252_));
  AND      g0236(.a(new_n88_), .b(i_2_6_111_0), .O(new_n253_));
  AND      g0237(.a(new_n217_), .b(new_n149_), .O(new_n254_));
  OR       g0238(.a(new_n254_), .b(new_n144_), .O(new_n255_));
  AND      g0239(.a(new_n255_), .b(new_n253_), .O(new_n256_));
  AND      g0240(.a(new_n19_), .b(i_2_6_32_0), .O(new_n257_));
  AND      g0241(.a(new_n257_), .b(new_n22_), .O(new_n258_));
  OR       g0242(.a(new_n258_), .b(new_n114_), .O(new_n259_));
  AND      g0243(.a(new_n259_), .b(new_n157_), .O(new_n260_));
  OR       g0244(.a(new_n144_), .b(new_n73_), .O(new_n261_));
  AND      g0245(.a(new_n261_), .b(i_2_6_32_0), .O(new_n262_));
  NOT      g0246(.a(new_n81_), .O(new_n263_));
  NAND     g0247(.a(new_n95_), .b(i_2_6_142_0), .O(new_n264_));
  NAND     g0248(.a(new_n264_), .b(new_n263_), .O(new_n265_));
  OR       g0249(.a(new_n265_), .b(new_n262_), .O(new_n266_));
  OR       g0250(.a(new_n266_), .b(new_n260_), .O(new_n267_));
  AND      g0251(.a(new_n267_), .b(i_2_6_34_0), .O(new_n268_));
  OR       g0252(.a(new_n268_), .b(new_n256_), .O(new_n269_));
  AND      g0253(.a(new_n269_), .b(new_n35_), .O(new_n270_));
  OR       g0254(.a(new_n270_), .b(new_n252_), .O(new_n271_));
  OR       g0255(.a(new_n22_), .b(i_2_6_40_0), .O(new_n272_));
  OR       g0256(.a(new_n272_), .b(i_2_6_142_0), .O(new_n273_));
  NAND     g0257(.a(new_n273_), .b(i_2_6_84_0), .O(new_n274_));
  AND      g0258(.a(new_n274_), .b(new_n214_), .O(new_n275_));
  OR       g0259(.a(i_2_6_124_0), .b(new_n22_), .O(new_n276_));
  OR       g0260(.a(new_n276_), .b(i_2_6_142_0), .O(new_n277_));
  OR       g0261(.a(new_n19_), .b(i_2_6_110_0), .O(new_n278_));
  AND      g0262(.a(new_n278_), .b(i_2_6_111_0), .O(new_n279_));
  AND      g0263(.a(new_n279_), .b(new_n277_), .O(new_n280_));
  OR       g0264(.a(new_n280_), .b(new_n275_), .O(new_n281_));
  AND      g0265(.a(new_n281_), .b(i_2_6_63_0), .O(new_n282_));
  AND      g0266(.a(new_n179_), .b(i_2_6_142_0), .O(new_n283_));
  OR       g0267(.a(new_n283_), .b(new_n282_), .O(new_n284_));
  AND      g0268(.a(new_n284_), .b(i_2_6_32_0), .O(new_n285_));
  NAND     g0269(.a(new_n195_), .b(new_n21_), .O(new_n286_));
  OR       g0270(.a(new_n28_), .b(i_2_6_110_0), .O(new_n287_));
  OR       g0271(.a(new_n287_), .b(new_n134_), .O(new_n288_));
  NAND     g0272(.a(new_n288_), .b(new_n286_), .O(new_n289_));
  AND      g0273(.a(new_n289_), .b(new_n22_), .O(new_n290_));
  AND      g0274(.a(new_n113_), .b(i_2_6_34_0), .O(new_n291_));
  OR       g0275(.a(new_n74_), .b(new_n36_), .O(new_n292_));
  AND      g0276(.a(new_n292_), .b(i_2_6_142_0), .O(new_n293_));
  OR       g0277(.a(new_n293_), .b(new_n291_), .O(new_n294_));
  OR       g0278(.a(new_n294_), .b(new_n290_), .O(new_n295_));
  OR       g0279(.a(new_n295_), .b(new_n285_), .O(new_n296_));
  AND      g0280(.a(new_n296_), .b(new_n18_), .O(new_n297_));
  OR       g0281(.a(new_n143_), .b(new_n47_), .O(new_n298_));
  AND      g0282(.a(new_n298_), .b(i_2_6_63_0), .O(new_n299_));
  OR       g0283(.a(i_2_6_124_0), .b(i_2_6_118_0), .O(new_n300_));
  NOT      g0284(.a(new_n300_), .O(new_n301_));
  OR       g0285(.a(new_n301_), .b(new_n178_), .O(new_n302_));
  AND      g0286(.a(new_n302_), .b(i_2_6_40_0), .O(new_n303_));
  OR       g0287(.a(new_n114_), .b(new_n95_), .O(new_n304_));
  OR       g0288(.a(new_n304_), .b(new_n303_), .O(new_n305_));
  NAND     g0289(.a(i_2_6_118_0), .b(i_2_6_84_0), .O(new_n306_));
  OR       g0290(.a(new_n306_), .b(new_n112_), .O(new_n307_));
  AND      g0291(.a(new_n307_), .b(new_n305_), .O(new_n308_));
  OR       g0292(.a(new_n68_), .b(new_n18_), .O(new_n309_));
  OR       g0293(.a(i_2_6_142_0), .b(i_2_6_110_0), .O(new_n310_));
  AND      g0294(.a(new_n310_), .b(new_n19_), .O(new_n311_));
  AND      g0295(.a(new_n311_), .b(new_n309_), .O(new_n312_));
  AND      g0296(.a(i_2_6_110_0), .b(i_2_6_32_0), .O(new_n313_));
  AND      g0297(.a(new_n313_), .b(new_n73_), .O(new_n314_));
  OR       g0298(.a(new_n314_), .b(new_n312_), .O(new_n315_));
  OR       g0299(.a(new_n315_), .b(new_n308_), .O(new_n316_));
  OR       g0300(.a(new_n316_), .b(new_n299_), .O(new_n317_));
  AND      g0301(.a(new_n317_), .b(i_2_6_62_0), .O(new_n318_));
  AND      g0302(.a(new_n19_), .b(i_2_6_111_0), .O(new_n319_));
  AND      g0303(.a(new_n319_), .b(i_2_6_110_0), .O(new_n320_));
  AND      g0304(.a(new_n320_), .b(new_n109_), .O(new_n321_));
  AND      g0305(.a(new_n310_), .b(new_n23_), .O(new_n322_));
  AND      g0306(.a(new_n322_), .b(new_n257_), .O(new_n323_));
  OR       g0307(.a(new_n323_), .b(new_n68_), .O(new_n324_));
  OR       g0308(.a(new_n324_), .b(new_n253_), .O(new_n325_));
  AND      g0309(.a(new_n325_), .b(i_2_6_63_0), .O(new_n326_));
  OR       g0310(.a(new_n326_), .b(new_n321_), .O(new_n327_));
  OR       g0311(.a(new_n327_), .b(new_n318_), .O(new_n328_));
  AND      g0312(.a(new_n328_), .b(i_2_6_34_0), .O(new_n329_));
  OR       g0313(.a(new_n329_), .b(new_n297_), .O(new_n330_));
  OR       g0314(.a(new_n330_), .b(new_n271_), .O(new_n331_));
  AND      g0315(.a(new_n331_), .b(i_2_6_33_0), .O(new_n332_));
  OR       g0316(.a(new_n332_), .b(new_n210_), .O(new_n333_));
  AND      g0317(.a(new_n333_), .b(new_n193_), .O(new_n334_));
  OR       g0318(.a(i_2_6_118_0), .b(i_2_6_84_0), .O(new_n335_));
  NOT      g0319(.a(new_n335_), .O(new_n336_));
  AND      g0320(.a(new_n19_), .b(i_2_6_110_0), .O(new_n337_));
  OR       g0321(.a(new_n337_), .b(i_2_6_111_0), .O(new_n338_));
  AND      g0322(.a(new_n338_), .b(new_n23_), .O(new_n339_));
  OR       g0323(.a(new_n339_), .b(i_2_6_111_0), .O(new_n340_));
  AND      g0324(.a(new_n340_), .b(i_2_6_142_0), .O(new_n341_));
  OR       g0325(.a(new_n149_), .b(new_n19_), .O(new_n342_));
  AND      g0326(.a(new_n342_), .b(new_n253_), .O(new_n343_));
  OR       g0327(.a(new_n343_), .b(new_n341_), .O(new_n344_));
  AND      g0328(.a(new_n344_), .b(i_2_6_32_0), .O(new_n345_));
  OR       g0329(.a(new_n345_), .b(new_n321_), .O(new_n346_));
  AND      g0330(.a(new_n346_), .b(i_2_6_62_0), .O(new_n347_));
  AND      g0331(.a(new_n85_), .b(new_n74_), .O(new_n348_));
  OR       g0332(.a(new_n348_), .b(new_n347_), .O(new_n349_));
  AND      g0333(.a(new_n349_), .b(new_n336_), .O(new_n350_));
  NAND     g0334(.a(new_n180_), .b(new_n27_), .O(new_n351_));
  AND      g0335(.a(new_n351_), .b(new_n18_), .O(new_n352_));
  OR       g0336(.a(new_n19_), .b(i_2_6_40_0), .O(new_n353_));
  OR       g0337(.a(i_2_6_142_0), .b(new_n18_), .O(new_n354_));
  OR       g0338(.a(new_n354_), .b(i_2_6_62_0), .O(new_n355_));
  OR       g0339(.a(new_n355_), .b(new_n353_), .O(new_n356_));
  NAND     g0340(.a(new_n356_), .b(new_n22_), .O(new_n357_));
  AND      g0341(.a(new_n357_), .b(new_n35_), .O(new_n358_));
  OR       g0342(.a(new_n358_), .b(new_n352_), .O(new_n359_));
  AND      g0343(.a(new_n359_), .b(i_2_6_32_0), .O(new_n360_));
  AND      g0344(.a(new_n18_), .b(i_2_6_62_0), .O(new_n361_));
  OR       g0345(.a(new_n310_), .b(i_2_6_84_0), .O(new_n362_));
  NOT      g0346(.a(new_n362_), .O(new_n363_));
  OR       g0347(.a(new_n363_), .b(new_n361_), .O(new_n364_));
  AND      g0348(.a(new_n364_), .b(i_2_6_32_0), .O(new_n365_));
  NOT      g0349(.a(new_n27_), .O(new_n366_));
  AND      g0350(.a(new_n247_), .b(new_n366_), .O(new_n367_));
  AND      g0351(.a(new_n81_), .b(new_n18_), .O(new_n368_));
  OR       g0352(.a(new_n368_), .b(new_n79_), .O(new_n369_));
  OR       g0353(.a(new_n369_), .b(new_n367_), .O(new_n370_));
  OR       g0354(.a(new_n370_), .b(new_n365_), .O(new_n371_));
  AND      g0355(.a(new_n371_), .b(new_n19_), .O(new_n372_));
  OR       g0356(.a(new_n361_), .b(i_2_6_84_0), .O(new_n373_));
  NAND     g0357(.a(new_n373_), .b(new_n164_), .O(new_n374_));
  AND      g0358(.a(new_n27_), .b(i_2_6_118_0), .O(new_n375_));
  OR       g0359(.a(new_n336_), .b(new_n73_), .O(new_n376_));
  NAND     g0360(.a(new_n376_), .b(i_2_6_110_0), .O(new_n377_));
  OR       g0361(.a(new_n377_), .b(new_n375_), .O(new_n378_));
  NAND     g0362(.a(new_n378_), .b(new_n374_), .O(new_n379_));
  OR       g0363(.a(new_n379_), .b(new_n372_), .O(new_n380_));
  OR       g0364(.a(new_n380_), .b(new_n360_), .O(new_n381_));
  AND      g0365(.a(new_n381_), .b(i_2_6_34_0), .O(new_n382_));
  OR       g0366(.a(new_n382_), .b(new_n350_), .O(new_n383_));
  AND      g0367(.a(new_n383_), .b(new_n193_), .O(new_n384_));
  AND      g0368(.a(new_n337_), .b(new_n58_), .O(new_n385_));
  OR       g0369(.a(i_2_6_84_0), .b(i_2_6_40_0), .O(new_n386_));
  NOT      g0370(.a(new_n386_), .O(new_n387_));
  AND      g0371(.a(new_n387_), .b(new_n385_), .O(new_n388_));
  OR       g0372(.a(new_n337_), .b(i_2_6_142_0), .O(new_n389_));
  AND      g0373(.a(new_n389_), .b(new_n166_), .O(new_n390_));
  OR       g0374(.a(new_n58_), .b(new_n35_), .O(new_n391_));
  AND      g0375(.a(new_n391_), .b(new_n149_), .O(new_n392_));
  AND      g0376(.a(new_n166_), .b(new_n50_), .O(new_n393_));
  OR       g0377(.a(new_n393_), .b(new_n392_), .O(new_n394_));
  OR       g0378(.a(new_n337_), .b(new_n35_), .O(new_n395_));
  OR       g0379(.a(new_n230_), .b(new_n179_), .O(new_n396_));
  AND      g0380(.a(new_n396_), .b(new_n395_), .O(new_n397_));
  AND      g0381(.a(new_n397_), .b(new_n151_), .O(new_n398_));
  AND      g0382(.a(new_n398_), .b(new_n394_), .O(new_n399_));
  OR       g0383(.a(new_n399_), .b(new_n390_), .O(new_n400_));
  AND      g0384(.a(new_n400_), .b(i_2_6_62_0), .O(new_n401_));
  OR       g0385(.a(new_n401_), .b(new_n388_), .O(new_n402_));
  AND      g0386(.a(new_n402_), .b(new_n18_), .O(new_n403_));
  OR       g0387(.a(new_n361_), .b(new_n149_), .O(new_n404_));
  AND      g0388(.a(new_n404_), .b(i_2_6_111_0), .O(new_n405_));
  OR       g0389(.a(i_2_6_111_0), .b(new_n20_), .O(new_n406_));
  OR       g0390(.a(new_n229_), .b(new_n26_), .O(new_n407_));
  NAND     g0391(.a(new_n407_), .b(new_n406_), .O(new_n408_));
  AND      g0392(.a(new_n408_), .b(new_n18_), .O(new_n409_));
  OR       g0393(.a(new_n409_), .b(new_n405_), .O(new_n410_));
  AND      g0394(.a(new_n410_), .b(new_n35_), .O(new_n411_));
  OR       g0395(.a(i_2_6_111_0), .b(i_2_6_84_0), .O(new_n412_));
  AND      g0396(.a(new_n19_), .b(i_2_6_62_0), .O(new_n413_));
  NAND     g0397(.a(new_n413_), .b(i_2_6_51_0), .O(new_n414_));
  AND      g0398(.a(new_n414_), .b(new_n412_), .O(new_n415_));
  OR       g0399(.a(new_n415_), .b(new_n20_), .O(new_n416_));
  AND      g0400(.a(new_n27_), .b(new_n19_), .O(new_n417_));
  OR       g0401(.a(new_n375_), .b(new_n23_), .O(new_n418_));
  OR       g0402(.a(new_n418_), .b(new_n417_), .O(new_n419_));
  NAND     g0403(.a(new_n419_), .b(new_n416_), .O(new_n420_));
  AND      g0404(.a(new_n420_), .b(i_2_6_142_0), .O(new_n421_));
  OR       g0405(.a(new_n413_), .b(new_n18_), .O(new_n422_));
  AND      g0406(.a(new_n342_), .b(i_2_6_111_0), .O(new_n423_));
  AND      g0407(.a(new_n423_), .b(new_n422_), .O(new_n424_));
  OR       g0408(.a(new_n424_), .b(new_n421_), .O(new_n425_));
  OR       g0409(.a(new_n425_), .b(new_n411_), .O(new_n426_));
  AND      g0410(.a(new_n426_), .b(i_2_6_32_0), .O(new_n427_));
  OR       g0411(.a(new_n427_), .b(new_n403_), .O(new_n428_));
  AND      g0412(.a(new_n428_), .b(i_2_6_34_0), .O(new_n429_));
  NOT      g0413(.a(new_n49_), .O(new_n430_));
  AND      g0414(.a(new_n361_), .b(new_n430_), .O(new_n431_));
  AND      g0415(.a(new_n431_), .b(new_n321_), .O(new_n432_));
  OR       g0416(.a(new_n432_), .b(new_n429_), .O(new_n433_));
  OR       g0417(.a(new_n433_), .b(new_n384_), .O(new_n434_));
  AND      g0418(.a(new_n434_), .b(i_2_6_63_0), .O(new_n435_));
  OR       g0419(.a(new_n435_), .b(new_n334_), .O(new_n436_));
  OR       g0420(.a(new_n436_), .b(new_n192_), .O(new_n437_));
  AND      g0421(.a(new_n437_), .b(i_2_6_5_0), .O(new_n438_));
  AND      g0422(.a(new_n94_), .b(i_2_6_110_0), .O(new_n439_));
  AND      g0423(.a(new_n140_), .b(i_2_6_111_0), .O(new_n440_));
  OR       g0424(.a(new_n440_), .b(new_n127_), .O(new_n441_));
  OR       g0425(.a(new_n441_), .b(new_n439_), .O(new_n442_));
  OR       g0426(.a(new_n442_), .b(new_n339_), .O(new_n443_));
  AND      g0427(.a(new_n443_), .b(i_2_6_32_0), .O(new_n444_));
  AND      g0428(.a(new_n149_), .b(i_2_6_142_0), .O(new_n445_));
  OR       g0429(.a(new_n445_), .b(new_n444_), .O(new_n446_));
  AND      g0430(.a(new_n446_), .b(i_2_6_63_0), .O(new_n447_));
  OR       g0431(.a(new_n447_), .b(new_n321_), .O(new_n448_));
  AND      g0432(.a(new_n448_), .b(new_n193_), .O(new_n449_));
  OR       g0433(.a(new_n74_), .b(new_n58_), .O(new_n450_));
  AND      g0434(.a(new_n450_), .b(new_n218_), .O(new_n451_));
  AND      g0435(.a(new_n18_), .b(i_2_6_63_0), .O(new_n452_));
  OR       g0436(.a(new_n322_), .b(new_n157_), .O(new_n453_));
  AND      g0437(.a(new_n453_), .b(new_n452_), .O(new_n454_));
  OR       g0438(.a(i_2_6_124_0), .b(i_2_6_51_0), .O(new_n455_));
  NOT      g0439(.a(new_n455_), .O(new_n456_));
  AND      g0440(.a(new_n456_), .b(i_2_6_40_0), .O(new_n457_));
  OR       g0441(.a(new_n457_), .b(new_n454_), .O(new_n458_));
  AND      g0442(.a(new_n458_), .b(new_n35_), .O(new_n459_));
  OR       g0443(.a(new_n459_), .b(new_n451_), .O(new_n460_));
  OR       g0444(.a(new_n460_), .b(new_n449_), .O(new_n461_));
  AND      g0445(.a(new_n461_), .b(i_2_6_33_0), .O(new_n462_));
  NOT      g0446(.a(i_2_6_5_0), .O(new_n463_));
  NOT      g0447(.a(new_n195_), .O(new_n464_));
  OR       g0448(.a(new_n56_), .b(new_n28_), .O(new_n465_));
  NAND     g0449(.a(new_n465_), .b(new_n464_), .O(new_n466_));
  AND      g0450(.a(new_n466_), .b(new_n463_), .O(new_n467_));
  OR       g0451(.a(i_2_6_110_0), .b(new_n193_), .O(new_n468_));
  OR       g0452(.a(new_n468_), .b(new_n272_), .O(new_n469_));
  NAND     g0453(.a(new_n56_), .b(i_2_6_33_0), .O(new_n470_));
  NAND     g0454(.a(new_n470_), .b(new_n469_), .O(new_n471_));
  OR       g0455(.a(new_n471_), .b(new_n467_), .O(new_n472_));
  AND      g0456(.a(new_n472_), .b(new_n19_), .O(new_n473_));
  OR       g0457(.a(i_2_6_111_0), .b(new_n193_), .O(new_n474_));
  AND      g0458(.a(new_n474_), .b(i_2_6_33_0), .O(new_n475_));
  AND      g0459(.a(new_n29_), .b(i_2_6_33_0), .O(new_n476_));
  AND      g0460(.a(new_n476_), .b(new_n24_), .O(new_n477_));
  OR       g0461(.a(new_n477_), .b(new_n475_), .O(new_n478_));
  OR       g0462(.a(new_n478_), .b(new_n473_), .O(new_n479_));
  AND      g0463(.a(new_n479_), .b(new_n18_), .O(new_n480_));
  OR       g0464(.a(new_n221_), .b(new_n22_), .O(new_n481_));
  OR       g0465(.a(i_2_6_124_0), .b(new_n20_), .O(new_n482_));
  AND      g0466(.a(new_n482_), .b(i_2_6_51_0), .O(new_n483_));
  AND      g0467(.a(new_n483_), .b(new_n481_), .O(new_n484_));
  AND      g0468(.a(new_n484_), .b(new_n58_), .O(new_n485_));
  AND      g0469(.a(new_n74_), .b(new_n18_), .O(new_n486_));
  OR       g0470(.a(new_n211_), .b(new_n19_), .O(new_n487_));
  OR       g0471(.a(i_2_6_111_0), .b(i_2_6_51_0), .O(new_n488_));
  NOT      g0472(.a(new_n488_), .O(new_n489_));
  AND      g0473(.a(new_n489_), .b(new_n487_), .O(new_n490_));
  AND      g0474(.a(i_2_6_142_0), .b(new_n22_), .O(new_n491_));
  OR       g0475(.a(i_2_6_51_0), .b(i_2_6_40_0), .O(new_n492_));
  NOT      g0476(.a(new_n492_), .O(new_n493_));
  OR       g0477(.a(new_n493_), .b(new_n491_), .O(new_n494_));
  AND      g0478(.a(new_n494_), .b(i_2_6_110_0), .O(new_n495_));
  OR       g0479(.a(new_n495_), .b(new_n490_), .O(new_n496_));
  OR       g0480(.a(new_n496_), .b(new_n486_), .O(new_n497_));
  OR       g0481(.a(new_n497_), .b(new_n485_), .O(new_n498_));
  AND      g0482(.a(new_n498_), .b(i_2_6_63_0), .O(new_n499_));
  OR       g0483(.a(new_n337_), .b(new_n193_), .O(new_n500_));
  OR       g0484(.a(new_n500_), .b(new_n279_), .O(new_n501_));
  OR       g0485(.a(new_n501_), .b(new_n151_), .O(new_n502_));
  AND      g0486(.a(new_n502_), .b(i_2_6_63_0), .O(new_n503_));
  OR       g0487(.a(new_n20_), .b(i_2_6_51_0), .O(new_n504_));
  OR       g0488(.a(new_n504_), .b(new_n28_), .O(new_n505_));
  AND      g0489(.a(new_n406_), .b(new_n322_), .O(new_n506_));
  AND      g0490(.a(i_2_6_111_0), .b(new_n193_), .O(new_n507_));
  OR       g0491(.a(new_n507_), .b(new_n68_), .O(new_n508_));
  NAND     g0492(.a(new_n508_), .b(new_n506_), .O(new_n509_));
  NAND     g0493(.a(new_n509_), .b(new_n505_), .O(new_n510_));
  OR       g0494(.a(new_n510_), .b(new_n503_), .O(new_n511_));
  AND      g0495(.a(new_n511_), .b(i_2_6_33_0), .O(new_n512_));
  OR       g0496(.a(new_n512_), .b(new_n499_), .O(new_n513_));
  OR       g0497(.a(new_n513_), .b(new_n480_), .O(new_n514_));
  AND      g0498(.a(new_n514_), .b(i_2_6_32_0), .O(new_n515_));
  NOT      g0499(.a(i_2_6_33_0), .O(new_n516_));
  OR       g0500(.a(new_n492_), .b(new_n516_), .O(new_n517_));
  AND      g0501(.a(i_2_6_142_0), .b(new_n193_), .O(new_n518_));
  OR       g0502(.a(new_n504_), .b(i_2_6_40_0), .O(new_n519_));
  NAND     g0503(.a(new_n519_), .b(new_n516_), .O(new_n520_));
  OR       g0504(.a(new_n310_), .b(new_n23_), .O(new_n521_));
  AND      g0505(.a(new_n521_), .b(new_n520_), .O(new_n522_));
  OR       g0506(.a(new_n522_), .b(new_n518_), .O(new_n523_));
  NAND     g0507(.a(new_n523_), .b(new_n18_), .O(new_n524_));
  NAND     g0508(.a(new_n524_), .b(new_n517_), .O(new_n525_));
  AND      g0509(.a(new_n525_), .b(i_2_6_63_0), .O(new_n526_));
  AND      g0510(.a(i_2_6_142_0), .b(i_2_6_33_0), .O(new_n527_));
  AND      g0511(.a(new_n527_), .b(new_n199_), .O(new_n528_));
  AND      g0512(.a(i_2_6_63_0), .b(i_2_6_33_0), .O(new_n529_));
  AND      g0513(.a(new_n529_), .b(new_n24_), .O(new_n530_));
  OR       g0514(.a(new_n144_), .b(i_2_6_33_0), .O(new_n531_));
  AND      g0515(.a(new_n531_), .b(new_n247_), .O(new_n532_));
  OR       g0516(.a(new_n532_), .b(new_n530_), .O(new_n533_));
  AND      g0517(.a(new_n533_), .b(i_2_6_110_0), .O(new_n534_));
  OR       g0518(.a(new_n504_), .b(new_n239_), .O(new_n535_));
  OR       g0519(.a(i_2_6_118_0), .b(new_n516_), .O(new_n536_));
  OR       g0520(.a(new_n536_), .b(new_n310_), .O(new_n537_));
  AND      g0521(.a(new_n537_), .b(new_n535_), .O(new_n538_));
  OR       g0522(.a(new_n538_), .b(new_n23_), .O(new_n539_));
  OR       g0523(.a(i_2_6_110_0), .b(i_2_6_32_0), .O(new_n540_));
  OR       g0524(.a(i_2_6_142_0), .b(i_2_6_51_0), .O(new_n541_));
  OR       g0525(.a(new_n541_), .b(new_n246_), .O(new_n542_));
  OR       g0526(.a(new_n542_), .b(new_n540_), .O(new_n543_));
  NAND     g0527(.a(new_n543_), .b(new_n539_), .O(new_n544_));
  OR       g0528(.a(new_n544_), .b(new_n534_), .O(new_n545_));
  AND      g0529(.a(new_n545_), .b(new_n19_), .O(new_n546_));
  OR       g0530(.a(new_n546_), .b(new_n528_), .O(new_n547_));
  OR       g0531(.a(new_n547_), .b(new_n526_), .O(new_n548_));
  AND      g0532(.a(new_n548_), .b(i_2_6_111_0), .O(new_n549_));
  OR       g0533(.a(new_n549_), .b(new_n515_), .O(new_n550_));
  AND      g0534(.a(new_n550_), .b(new_n35_), .O(new_n551_));
  NAND     g0535(.a(new_n103_), .b(i_2_6_142_0), .O(new_n552_));
  NAND     g0536(.a(new_n541_), .b(i_2_6_40_0), .O(new_n553_));
  NAND     g0537(.a(new_n553_), .b(new_n476_), .O(new_n554_));
  NAND     g0538(.a(new_n554_), .b(new_n552_), .O(new_n555_));
  AND      g0539(.a(new_n555_), .b(i_2_6_110_0), .O(new_n556_));
  AND      g0540(.a(i_2_6_111_0), .b(i_2_6_33_0), .O(new_n557_));
  AND      g0541(.a(new_n557_), .b(new_n493_), .O(new_n558_));
  OR       g0542(.a(new_n507_), .b(i_2_6_33_0), .O(new_n559_));
  AND      g0543(.a(new_n559_), .b(new_n109_), .O(new_n560_));
  OR       g0544(.a(new_n560_), .b(new_n475_), .O(new_n561_));
  AND      g0545(.a(new_n561_), .b(i_2_6_63_0), .O(new_n562_));
  OR       g0546(.a(new_n562_), .b(new_n558_), .O(new_n563_));
  OR       g0547(.a(new_n563_), .b(new_n556_), .O(new_n564_));
  AND      g0548(.a(new_n564_), .b(new_n19_), .O(new_n565_));
  AND      g0549(.a(new_n475_), .b(new_n144_), .O(new_n566_));
  NOT      g0550(.a(new_n504_), .O(new_n567_));
  NOT      g0551(.a(new_n72_), .O(new_n568_));
  OR       g0552(.a(new_n234_), .b(new_n28_), .O(new_n569_));
  NAND     g0553(.a(new_n569_), .b(new_n568_), .O(new_n570_));
  AND      g0554(.a(new_n570_), .b(new_n567_), .O(new_n571_));
  OR       g0555(.a(new_n58_), .b(i_2_6_63_0), .O(new_n572_));
  AND      g0556(.a(new_n572_), .b(new_n193_), .O(new_n573_));
  AND      g0557(.a(new_n69_), .b(i_2_6_111_0), .O(new_n574_));
  OR       g0558(.a(new_n574_), .b(new_n573_), .O(new_n575_));
  AND      g0559(.a(new_n575_), .b(i_2_6_33_0), .O(new_n576_));
  OR       g0560(.a(new_n576_), .b(new_n571_), .O(new_n577_));
  AND      g0561(.a(new_n577_), .b(new_n23_), .O(new_n578_));
  OR       g0562(.a(new_n578_), .b(new_n566_), .O(new_n579_));
  OR       g0563(.a(new_n579_), .b(new_n565_), .O(new_n580_));
  AND      g0564(.a(new_n580_), .b(i_2_6_32_0), .O(new_n581_));
  AND      g0565(.a(new_n81_), .b(new_n193_), .O(new_n582_));
  AND      g0566(.a(new_n582_), .b(new_n527_), .O(new_n583_));
  AND      g0567(.a(new_n22_), .b(i_2_6_110_0), .O(new_n584_));
  AND      g0568(.a(new_n493_), .b(new_n127_), .O(new_n585_));
  AND      g0569(.a(new_n585_), .b(new_n584_), .O(new_n586_));
  AND      g0570(.a(new_n310_), .b(new_n319_), .O(new_n587_));
  NOT      g0571(.a(new_n68_), .O(new_n588_));
  AND      g0572(.a(new_n588_), .b(i_2_6_40_0), .O(new_n589_));
  NOT      g0573(.a(new_n589_), .O(new_n590_));
  AND      g0574(.a(new_n590_), .b(new_n587_), .O(new_n591_));
  OR       g0575(.a(new_n585_), .b(new_n507_), .O(new_n592_));
  OR       g0576(.a(new_n592_), .b(new_n591_), .O(new_n593_));
  AND      g0577(.a(new_n593_), .b(i_2_6_33_0), .O(new_n594_));
  OR       g0578(.a(new_n594_), .b(new_n586_), .O(new_n595_));
  AND      g0579(.a(new_n595_), .b(i_2_6_63_0), .O(new_n596_));
  OR       g0580(.a(new_n596_), .b(new_n583_), .O(new_n597_));
  OR       g0581(.a(new_n597_), .b(new_n581_), .O(new_n598_));
  AND      g0582(.a(new_n598_), .b(new_n18_), .O(new_n599_));
  OR       g0583(.a(new_n599_), .b(new_n551_), .O(new_n600_));
  OR       g0584(.a(new_n600_), .b(new_n462_), .O(new_n601_));
  AND      g0585(.a(new_n601_), .b(i_2_6_34_0), .O(new_n602_));
  NAND     g0586(.a(new_n149_), .b(i_2_6_124_0), .O(new_n603_));
  OR       g0587(.a(new_n603_), .b(i_2_6_5_0), .O(new_n604_));
  AND      g0588(.a(new_n88_), .b(i_2_6_32_0), .O(new_n605_));
  NAND     g0589(.a(new_n605_), .b(new_n456_), .O(new_n606_));
  NAND     g0590(.a(new_n606_), .b(new_n604_), .O(new_n607_));
  NOT      g0591(.a(new_n536_), .O(new_n608_));
  AND      g0592(.a(new_n608_), .b(new_n59_), .O(new_n609_));
  AND      g0593(.a(new_n609_), .b(new_n607_), .O(new_n610_));
  AND      g0594(.a(new_n88_), .b(new_n18_), .O(new_n611_));
  NAND     g0595(.a(new_n112_), .b(new_n193_), .O(new_n612_));
  NOT      g0596(.a(new_n612_), .O(new_n613_));
  AND      g0597(.a(new_n613_), .b(new_n611_), .O(new_n614_));
  AND      g0598(.a(new_n69_), .b(new_n193_), .O(new_n615_));
  OR       g0599(.a(new_n615_), .b(new_n144_), .O(new_n616_));
  AND      g0600(.a(new_n616_), .b(new_n194_), .O(new_n617_));
  AND      g0601(.a(i_2_6_63_0), .b(new_n193_), .O(new_n618_));
  NAND     g0602(.a(new_n618_), .b(i_2_6_142_0), .O(new_n619_));
  OR       g0603(.a(new_n619_), .b(i_2_6_110_0), .O(new_n620_));
  AND      g0604(.a(new_n535_), .b(i_2_6_32_0), .O(new_n621_));
  AND      g0605(.a(new_n287_), .b(new_n21_), .O(new_n622_));
  OR       g0606(.a(new_n622_), .b(i_2_6_40_0), .O(new_n623_));
  OR       g0607(.a(new_n623_), .b(new_n621_), .O(new_n624_));
  NAND     g0608(.a(new_n624_), .b(new_n620_), .O(new_n625_));
  OR       g0609(.a(new_n625_), .b(new_n617_), .O(new_n626_));
  AND      g0610(.a(new_n626_), .b(new_n19_), .O(new_n627_));
  OR       g0611(.a(new_n627_), .b(new_n614_), .O(new_n628_));
  AND      g0612(.a(new_n628_), .b(i_2_6_111_0), .O(new_n629_));
  NOT      g0613(.a(new_n619_), .O(new_n630_));
  OR       g0614(.a(new_n18_), .b(i_2_6_110_0), .O(new_n631_));
  NAND     g0615(.a(new_n631_), .b(new_n257_), .O(new_n632_));
  NAND     g0616(.a(new_n632_), .b(new_n603_), .O(new_n633_));
  AND      g0617(.a(new_n633_), .b(new_n630_), .O(new_n634_));
  OR       g0618(.a(new_n634_), .b(new_n629_), .O(new_n635_));
  AND      g0619(.a(new_n35_), .b(i_2_6_33_0), .O(new_n636_));
  AND      g0620(.a(new_n636_), .b(new_n635_), .O(new_n637_));
  OR       g0621(.a(new_n637_), .b(new_n610_), .O(new_n638_));
  OR       g0622(.a(new_n638_), .b(new_n602_), .O(new_n639_));
  AND      g0623(.a(new_n639_), .b(i_2_6_62_0), .O(new_n640_));
  AND      g0624(.a(new_n337_), .b(new_n18_), .O(new_n641_));
  AND      g0625(.a(new_n641_), .b(new_n493_), .O(new_n642_));
  AND      g0626(.a(new_n642_), .b(i_2_6_142_0), .O(new_n643_));
  NAND     g0627(.a(new_n194_), .b(new_n193_), .O(new_n644_));
  OR       g0628(.a(new_n127_), .b(new_n23_), .O(new_n645_));
  AND      g0629(.a(new_n645_), .b(new_n194_), .O(new_n646_));
  OR       g0630(.a(new_n646_), .b(new_n585_), .O(new_n647_));
  NAND     g0631(.a(new_n647_), .b(i_2_6_110_0), .O(new_n648_));
  NAND     g0632(.a(new_n648_), .b(new_n644_), .O(new_n649_));
  AND      g0633(.a(new_n649_), .b(new_n35_), .O(new_n650_));
  OR       g0634(.a(new_n650_), .b(new_n643_), .O(new_n651_));
  AND      g0635(.a(new_n651_), .b(i_2_6_111_0), .O(new_n652_));
  AND      g0636(.a(new_n591_), .b(new_n336_), .O(new_n653_));
  OR       g0637(.a(new_n46_), .b(new_n18_), .O(new_n654_));
  AND      g0638(.a(new_n654_), .b(new_n319_), .O(new_n655_));
  OR       g0639(.a(new_n179_), .b(new_n135_), .O(new_n656_));
  OR       g0640(.a(new_n247_), .b(new_n73_), .O(new_n657_));
  AND      g0641(.a(new_n657_), .b(new_n656_), .O(new_n658_));
  OR       g0642(.a(new_n658_), .b(new_n655_), .O(new_n659_));
  AND      g0643(.a(new_n659_), .b(i_2_6_142_0), .O(new_n660_));
  AND      g0644(.a(new_n376_), .b(new_n46_), .O(new_n661_));
  OR       g0645(.a(new_n661_), .b(new_n368_), .O(new_n662_));
  OR       g0646(.a(new_n662_), .b(new_n660_), .O(new_n663_));
  AND      g0647(.a(new_n663_), .b(i_2_6_32_0), .O(new_n664_));
  OR       g0648(.a(new_n664_), .b(new_n653_), .O(new_n665_));
  AND      g0649(.a(new_n665_), .b(i_2_6_63_0), .O(new_n666_));
  OR       g0650(.a(new_n666_), .b(new_n652_), .O(new_n667_));
  AND      g0651(.a(new_n667_), .b(i_2_6_34_0), .O(new_n668_));
  OR       g0652(.a(new_n387_), .b(new_n81_), .O(new_n669_));
  AND      g0653(.a(new_n669_), .b(new_n40_), .O(new_n670_));
  AND      g0654(.a(new_n195_), .b(new_n22_), .O(new_n671_));
  OR       g0655(.a(new_n671_), .b(new_n166_), .O(new_n672_));
  AND      g0656(.a(new_n672_), .b(new_n18_), .O(new_n673_));
  OR       g0657(.a(new_n673_), .b(new_n670_), .O(new_n674_));
  AND      g0658(.a(new_n674_), .b(new_n19_), .O(new_n675_));
  NOT      g0659(.a(new_n88_), .O(new_n676_));
  AND      g0660(.a(new_n676_), .b(i_2_6_34_0), .O(new_n677_));
  AND      g0661(.a(new_n677_), .b(new_n160_), .O(new_n678_));
  OR       g0662(.a(new_n678_), .b(new_n675_), .O(new_n679_));
  AND      g0663(.a(new_n679_), .b(i_2_6_142_0), .O(new_n680_));
  AND      g0664(.a(new_n306_), .b(i_2_6_32_0), .O(new_n681_));
  OR       g0665(.a(new_n681_), .b(new_n397_), .O(new_n682_));
  AND      g0666(.a(new_n682_), .b(i_2_6_111_0), .O(new_n683_));
  AND      g0667(.a(new_n395_), .b(new_n247_), .O(new_n684_));
  OR       g0668(.a(new_n684_), .b(new_n683_), .O(new_n685_));
  AND      g0669(.a(new_n685_), .b(i_2_6_34_0), .O(new_n686_));
  NAND     g0670(.a(new_n412_), .b(new_n273_), .O(new_n687_));
  AND      g0671(.a(new_n687_), .b(i_2_6_32_0), .O(new_n688_));
  OR       g0672(.a(new_n688_), .b(new_n158_), .O(new_n689_));
  AND      g0673(.a(new_n689_), .b(new_n641_), .O(new_n690_));
  OR       g0674(.a(new_n690_), .b(new_n686_), .O(new_n691_));
  OR       g0675(.a(new_n691_), .b(new_n680_), .O(new_n692_));
  AND      g0676(.a(new_n692_), .b(new_n193_), .O(new_n693_));
  AND      g0677(.a(new_n28_), .b(i_2_6_110_0), .O(new_n694_));
  AND      g0678(.a(new_n301_), .b(new_n694_), .O(new_n695_));
  AND      g0679(.a(new_n695_), .b(new_n149_), .O(new_n696_));
  AND      g0680(.a(new_n696_), .b(new_n167_), .O(new_n697_));
  OR       g0681(.a(new_n697_), .b(new_n693_), .O(new_n698_));
  AND      g0682(.a(new_n698_), .b(i_2_6_63_0), .O(new_n699_));
  OR       g0683(.a(new_n699_), .b(new_n668_), .O(new_n700_));
  AND      g0684(.a(new_n700_), .b(i_2_6_33_0), .O(new_n701_));
  AND      g0685(.a(new_n688_), .b(i_2_6_124_0), .O(new_n702_));
  NAND     g0686(.a(new_n264_), .b(new_n21_), .O(new_n703_));
  AND      g0687(.a(new_n703_), .b(new_n35_), .O(new_n704_));
  OR       g0688(.a(new_n704_), .b(new_n702_), .O(new_n705_));
  AND      g0689(.a(new_n705_), .b(new_n18_), .O(new_n706_));
  AND      g0690(.a(new_n211_), .b(new_n22_), .O(new_n707_));
  AND      g0691(.a(new_n707_), .b(new_n136_), .O(new_n708_));
  OR       g0692(.a(new_n708_), .b(new_n706_), .O(new_n709_));
  AND      g0693(.a(new_n709_), .b(i_2_6_110_0), .O(new_n710_));
  AND      g0694(.a(new_n37_), .b(new_n18_), .O(new_n711_));
  OR       g0695(.a(new_n711_), .b(new_n710_), .O(new_n712_));
  AND      g0696(.a(new_n193_), .b(i_2_6_34_0), .O(new_n713_));
  AND      g0697(.a(new_n713_), .b(new_n712_), .O(new_n714_));
  OR       g0698(.a(new_n714_), .b(new_n701_), .O(new_n715_));
  OR       g0699(.a(new_n715_), .b(new_n640_), .O(new_n716_));
  OR       g0700(.a(new_n716_), .b(new_n438_), .O(new_n717_));
  AND      g0701(.a(new_n717_), .b(new_n17_), .O(new_n718_));
  NAND     g0702(.a(i_2_6_40_0), .b(i_2_6_5_0), .O(new_n719_));
  NAND     g0703(.a(new_n719_), .b(i_2_6_118_0), .O(new_n720_));
  AND      g0704(.a(new_n720_), .b(new_n319_), .O(new_n721_));
  AND      g0705(.a(new_n73_), .b(i_2_6_5_0), .O(new_n722_));
  OR       g0706(.a(i_2_6_118_0), .b(new_n463_), .O(new_n723_));
  NAND     g0707(.a(new_n723_), .b(new_n272_), .O(new_n724_));
  AND      g0708(.a(new_n724_), .b(i_2_6_142_0), .O(new_n725_));
  OR       g0709(.a(new_n725_), .b(new_n722_), .O(new_n726_));
  OR       g0710(.a(new_n726_), .b(new_n721_), .O(new_n727_));
  AND      g0711(.a(new_n727_), .b(i_2_6_110_0), .O(new_n728_));
  NAND     g0712(.a(new_n504_), .b(new_n300_), .O(new_n729_));
  AND      g0713(.a(new_n729_), .b(i_2_6_5_0), .O(new_n730_));
  OR       g0714(.a(new_n730_), .b(new_n368_), .O(new_n731_));
  AND      g0715(.a(new_n731_), .b(new_n24_), .O(new_n732_));
  AND      g0716(.a(i_2_6_110_0), .b(i_2_6_5_0), .O(new_n733_));
  OR       g0717(.a(new_n733_), .b(new_n440_), .O(new_n734_));
  AND      g0718(.a(new_n734_), .b(new_n247_), .O(new_n735_));
  OR       g0719(.a(new_n17_), .b(i_2_6_40_0), .O(new_n736_));
  OR       g0720(.a(new_n736_), .b(new_n28_), .O(new_n737_));
  NAND     g0721(.a(new_n737_), .b(new_n723_), .O(new_n738_));
  AND      g0722(.a(new_n738_), .b(new_n500_), .O(new_n739_));
  OR       g0723(.a(new_n733_), .b(new_n58_), .O(new_n740_));
  AND      g0724(.a(new_n740_), .b(new_n456_), .O(new_n741_));
  OR       g0725(.a(new_n741_), .b(new_n739_), .O(new_n742_));
  OR       g0726(.a(new_n742_), .b(new_n735_), .O(new_n743_));
  OR       g0727(.a(new_n743_), .b(new_n732_), .O(new_n744_));
  OR       g0728(.a(new_n744_), .b(new_n728_), .O(new_n745_));
  AND      g0729(.a(new_n745_), .b(i_2_6_63_0), .O(new_n746_));
  AND      g0730(.a(new_n507_), .b(i_2_6_5_0), .O(new_n747_));
  AND      g0731(.a(new_n24_), .b(new_n193_), .O(new_n748_));
  OR       g0732(.a(new_n748_), .b(new_n18_), .O(new_n749_));
  OR       g0733(.a(new_n749_), .b(new_n109_), .O(new_n750_));
  AND      g0734(.a(new_n750_), .b(i_2_6_5_0), .O(new_n751_));
  AND      g0735(.a(new_n749_), .b(i_2_6_111_0), .O(new_n752_));
  OR       g0736(.a(new_n752_), .b(new_n751_), .O(new_n753_));
  AND      g0737(.a(new_n753_), .b(i_2_6_63_0), .O(new_n754_));
  OR       g0738(.a(new_n754_), .b(new_n747_), .O(new_n755_));
  AND      g0739(.a(new_n755_), .b(i_2_6_32_0), .O(new_n756_));
  AND      g0740(.a(i_2_6_124_0), .b(new_n193_), .O(new_n757_));
  OR       g0741(.a(new_n757_), .b(i_2_6_5_0), .O(new_n758_));
  AND      g0742(.a(new_n758_), .b(i_2_6_111_0), .O(new_n759_));
  AND      g0743(.a(new_n567_), .b(i_2_6_142_0), .O(new_n760_));
  OR       g0744(.a(new_n585_), .b(new_n760_), .O(new_n761_));
  OR       g0745(.a(new_n761_), .b(new_n759_), .O(new_n762_));
  AND      g0746(.a(new_n762_), .b(new_n18_), .O(new_n763_));
  OR       g0747(.a(new_n763_), .b(new_n756_), .O(new_n764_));
  OR       g0748(.a(new_n764_), .b(new_n746_), .O(new_n765_));
  AND      g0749(.a(new_n765_), .b(i_2_6_33_0), .O(new_n766_));
  NOT      g0750(.a(new_n736_), .O(new_n767_));
  OR       g0751(.a(new_n767_), .b(new_n475_), .O(new_n768_));
  AND      g0752(.a(new_n768_), .b(i_2_6_63_0), .O(new_n769_));
  AND      g0753(.a(new_n720_), .b(i_2_6_33_0), .O(new_n770_));
  OR       g0754(.a(new_n770_), .b(new_n20_), .O(new_n771_));
  OR       g0755(.a(new_n771_), .b(new_n769_), .O(new_n772_));
  OR       g0756(.a(i_2_6_51_0), .b(i_2_6_33_0), .O(new_n773_));
  OR       g0757(.a(i_2_6_118_0), .b(new_n239_), .O(new_n774_));
  OR       g0758(.a(new_n17_), .b(i_2_6_111_0), .O(new_n775_));
  OR       g0759(.a(new_n775_), .b(new_n774_), .O(new_n776_));
  NAND     g0760(.a(new_n776_), .b(new_n773_), .O(new_n777_));
  AND      g0761(.a(new_n777_), .b(new_n463_), .O(new_n778_));
  OR       g0762(.a(new_n778_), .b(i_2_6_110_0), .O(new_n779_));
  AND      g0763(.a(new_n779_), .b(i_2_6_142_0), .O(new_n780_));
  AND      g0764(.a(new_n780_), .b(new_n772_), .O(new_n781_));
  NAND     g0765(.a(new_n541_), .b(new_n66_), .O(new_n782_));
  AND      g0766(.a(new_n782_), .b(new_n23_), .O(new_n783_));
  OR       g0767(.a(new_n783_), .b(new_n618_), .O(new_n784_));
  AND      g0768(.a(new_n784_), .b(i_2_6_33_0), .O(new_n785_));
  OR       g0769(.a(new_n736_), .b(new_n310_), .O(new_n786_));
  NAND     g0770(.a(new_n786_), .b(new_n463_), .O(new_n787_));
  OR       g0771(.a(new_n452_), .b(new_n20_), .O(new_n788_));
  AND      g0772(.a(new_n788_), .b(i_2_6_5_0), .O(new_n789_));
  OR       g0773(.a(new_n789_), .b(new_n193_), .O(new_n790_));
  AND      g0774(.a(new_n790_), .b(new_n787_), .O(new_n791_));
  OR       g0775(.a(new_n791_), .b(new_n785_), .O(new_n792_));
  AND      g0776(.a(new_n792_), .b(i_2_6_111_0), .O(new_n793_));
  AND      g0777(.a(new_n468_), .b(i_2_6_5_0), .O(new_n794_));
  OR       g0778(.a(new_n794_), .b(new_n611_), .O(new_n795_));
  AND      g0779(.a(new_n795_), .b(i_2_6_33_0), .O(new_n796_));
  AND      g0780(.a(new_n567_), .b(new_n18_), .O(new_n797_));
  OR       g0781(.a(new_n797_), .b(new_n796_), .O(new_n798_));
  AND      g0782(.a(new_n798_), .b(i_2_6_63_0), .O(new_n799_));
  OR       g0783(.a(new_n799_), .b(new_n793_), .O(new_n800_));
  OR       g0784(.a(new_n800_), .b(new_n781_), .O(new_n801_));
  AND      g0785(.a(new_n801_), .b(new_n19_), .O(new_n802_));
  OR       g0786(.a(new_n529_), .b(new_n58_), .O(new_n803_));
  AND      g0787(.a(new_n803_), .b(new_n23_), .O(new_n804_));
  OR       g0788(.a(new_n475_), .b(new_n182_), .O(new_n805_));
  AND      g0789(.a(new_n805_), .b(i_2_6_63_0), .O(new_n806_));
  OR       g0790(.a(new_n806_), .b(new_n804_), .O(new_n807_));
  AND      g0791(.a(new_n807_), .b(i_2_6_5_0), .O(new_n808_));
  AND      g0792(.a(new_n618_), .b(new_n58_), .O(new_n809_));
  AND      g0793(.a(new_n809_), .b(new_n18_), .O(new_n810_));
  OR       g0794(.a(new_n72_), .b(new_n18_), .O(new_n811_));
  NAND     g0795(.a(new_n811_), .b(new_n193_), .O(new_n812_));
  AND      g0796(.a(new_n774_), .b(i_2_6_40_0), .O(new_n813_));
  OR       g0797(.a(new_n507_), .b(new_n18_), .O(new_n814_));
  NAND     g0798(.a(new_n814_), .b(i_2_6_142_0), .O(new_n815_));
  OR       g0799(.a(new_n815_), .b(new_n813_), .O(new_n816_));
  NAND     g0800(.a(new_n816_), .b(new_n812_), .O(new_n817_));
  AND      g0801(.a(new_n817_), .b(i_2_6_33_0), .O(new_n818_));
  OR       g0802(.a(new_n818_), .b(new_n810_), .O(new_n819_));
  OR       g0803(.a(new_n819_), .b(new_n808_), .O(new_n820_));
  AND      g0804(.a(new_n820_), .b(i_2_6_110_0), .O(new_n821_));
  OR       g0805(.a(new_n821_), .b(new_n802_), .O(new_n822_));
  AND      g0806(.a(new_n822_), .b(i_2_6_32_0), .O(new_n823_));
  OR       g0807(.a(i_2_6_118_0), .b(i_2_6_51_0), .O(new_n824_));
  NOT      g0808(.a(new_n824_), .O(new_n825_));
  OR       g0809(.a(new_n825_), .b(new_n254_), .O(new_n826_));
  AND      g0810(.a(new_n826_), .b(new_n58_), .O(new_n827_));
  AND      g0811(.a(new_n493_), .b(i_2_6_33_0), .O(new_n828_));
  AND      g0812(.a(new_n828_), .b(new_n278_), .O(new_n829_));
  AND      g0813(.a(new_n829_), .b(new_n389_), .O(new_n830_));
  OR       g0814(.a(new_n830_), .b(new_n827_), .O(new_n831_));
  AND      g0815(.a(new_n831_), .b(i_2_6_5_0), .O(new_n832_));
  OR       g0816(.a(new_n832_), .b(new_n823_), .O(new_n833_));
  OR       g0817(.a(new_n833_), .b(new_n766_), .O(new_n834_));
  AND      g0818(.a(new_n834_), .b(new_n35_), .O(new_n835_));
  NAND     g0819(.a(i_2_6_32_0), .b(i_2_6_5_0), .O(new_n836_));
  NOT      g0820(.a(new_n836_), .O(new_n837_));
  AND      g0821(.a(new_n837_), .b(new_n78_), .O(new_n838_));
  AND      g0822(.a(new_n507_), .b(new_n18_), .O(new_n839_));
  OR       g0823(.a(new_n839_), .b(new_n838_), .O(new_n840_));
  AND      g0824(.a(new_n840_), .b(i_2_6_40_0), .O(new_n841_));
  OR       g0825(.a(new_n199_), .b(new_n193_), .O(new_n842_));
  AND      g0826(.a(new_n842_), .b(i_2_6_5_0), .O(new_n843_));
  OR       g0827(.a(new_n194_), .b(new_n193_), .O(new_n844_));
  AND      g0828(.a(new_n844_), .b(i_2_6_111_0), .O(new_n845_));
  OR       g0829(.a(new_n845_), .b(new_n843_), .O(new_n846_));
  AND      g0830(.a(new_n846_), .b(new_n23_), .O(new_n847_));
  AND      g0831(.a(new_n474_), .b(i_2_6_110_0), .O(new_n848_));
  AND      g0832(.a(new_n814_), .b(i_2_6_32_0), .O(new_n849_));
  AND      g0833(.a(new_n849_), .b(new_n848_), .O(new_n850_));
  OR       g0834(.a(new_n850_), .b(new_n847_), .O(new_n851_));
  AND      g0835(.a(new_n851_), .b(i_2_6_63_0), .O(new_n852_));
  OR       g0836(.a(new_n852_), .b(new_n841_), .O(new_n853_));
  AND      g0837(.a(new_n853_), .b(new_n19_), .O(new_n854_));
  OR       g0838(.a(new_n582_), .b(new_n452_), .O(new_n855_));
  AND      g0839(.a(new_n855_), .b(i_2_6_32_0), .O(new_n856_));
  OR       g0840(.a(new_n848_), .b(new_n825_), .O(new_n857_));
  AND      g0841(.a(new_n857_), .b(i_2_6_63_0), .O(new_n858_));
  OR       g0842(.a(new_n858_), .b(new_n856_), .O(new_n859_));
  AND      g0843(.a(new_n859_), .b(i_2_6_5_0), .O(new_n860_));
  OR       g0844(.a(new_n112_), .b(new_n18_), .O(new_n861_));
  AND      g0845(.a(new_n861_), .b(new_n582_), .O(new_n862_));
  OR       g0846(.a(new_n862_), .b(new_n860_), .O(new_n863_));
  AND      g0847(.a(new_n863_), .b(new_n23_), .O(new_n864_));
  NAND     g0848(.a(new_n540_), .b(i_2_6_5_0), .O(new_n865_));
  NAND     g0849(.a(new_n865_), .b(new_n612_), .O(new_n866_));
  AND      g0850(.a(new_n866_), .b(i_2_6_111_0), .O(new_n867_));
  AND      g0851(.a(new_n733_), .b(new_n618_), .O(new_n868_));
  OR       g0852(.a(new_n868_), .b(new_n867_), .O(new_n869_));
  AND      g0853(.a(new_n869_), .b(new_n18_), .O(new_n870_));
  OR       g0854(.a(new_n870_), .b(new_n864_), .O(new_n871_));
  OR       g0855(.a(new_n871_), .b(new_n854_), .O(new_n872_));
  AND      g0856(.a(new_n872_), .b(i_2_6_142_0), .O(new_n873_));
  OR       g0857(.a(new_n618_), .b(new_n206_), .O(new_n874_));
  AND      g0858(.a(new_n874_), .b(new_n605_), .O(new_n875_));
  AND      g0859(.a(new_n468_), .b(new_n19_), .O(new_n876_));
  AND      g0860(.a(new_n876_), .b(new_n788_), .O(new_n877_));
  OR       g0861(.a(new_n877_), .b(new_n875_), .O(new_n878_));
  AND      g0862(.a(new_n878_), .b(i_2_6_111_0), .O(new_n879_));
  NAND     g0863(.a(new_n644_), .b(i_2_6_124_0), .O(new_n880_));
  OR       g0864(.a(new_n567_), .b(new_n194_), .O(new_n881_));
  AND      g0865(.a(new_n881_), .b(new_n95_), .O(new_n882_));
  AND      g0866(.a(new_n882_), .b(new_n880_), .O(new_n883_));
  OR       g0867(.a(new_n883_), .b(new_n879_), .O(new_n884_));
  AND      g0868(.a(new_n884_), .b(i_2_6_5_0), .O(new_n885_));
  AND      g0869(.a(new_n767_), .b(new_n695_), .O(new_n886_));
  OR       g0870(.a(new_n611_), .b(new_n19_), .O(new_n887_));
  OR       g0871(.a(new_n149_), .b(new_n18_), .O(new_n888_));
  AND      g0872(.a(new_n888_), .b(new_n618_), .O(new_n889_));
  AND      g0873(.a(new_n889_), .b(new_n887_), .O(new_n890_));
  OR       g0874(.a(new_n890_), .b(new_n886_), .O(new_n891_));
  AND      g0875(.a(new_n891_), .b(i_2_6_32_0), .O(new_n892_));
  OR       g0876(.a(new_n892_), .b(new_n642_), .O(new_n893_));
  AND      g0877(.a(new_n893_), .b(i_2_6_111_0), .O(new_n894_));
  OR       g0878(.a(new_n894_), .b(new_n885_), .O(new_n895_));
  OR       g0879(.a(new_n895_), .b(new_n873_), .O(new_n896_));
  AND      g0880(.a(new_n896_), .b(i_2_6_33_0), .O(new_n897_));
  AND      g0881(.a(new_n81_), .b(i_2_6_120_0), .O(new_n898_));
  AND      g0882(.a(new_n898_), .b(new_n643_), .O(new_n899_));
  NAND     g0883(.a(new_n236_), .b(new_n20_), .O(new_n900_));
  AND      g0884(.a(new_n825_), .b(i_2_6_142_0), .O(new_n901_));
  AND      g0885(.a(new_n901_), .b(new_n900_), .O(new_n902_));
  AND      g0886(.a(new_n572_), .b(i_2_6_118_0), .O(new_n903_));
  AND      g0887(.a(new_n903_), .b(new_n587_), .O(new_n904_));
  OR       g0888(.a(new_n904_), .b(new_n902_), .O(new_n905_));
  AND      g0889(.a(new_n905_), .b(new_n23_), .O(new_n906_));
  AND      g0890(.a(new_n103_), .b(i_2_6_142_0), .O(new_n907_));
  OR       g0891(.a(new_n907_), .b(new_n320_), .O(new_n908_));
  AND      g0892(.a(new_n908_), .b(new_n193_), .O(new_n909_));
  AND      g0893(.a(i_2_6_124_0), .b(i_2_6_120_0), .O(new_n910_));
  AND      g0894(.a(new_n910_), .b(new_n584_), .O(new_n911_));
  AND      g0895(.a(new_n911_), .b(new_n144_), .O(new_n912_));
  OR       g0896(.a(new_n912_), .b(new_n909_), .O(new_n913_));
  AND      g0897(.a(new_n913_), .b(new_n18_), .O(new_n914_));
  OR       g0898(.a(new_n914_), .b(new_n809_), .O(new_n915_));
  OR       g0899(.a(new_n915_), .b(new_n906_), .O(new_n916_));
  AND      g0900(.a(new_n916_), .b(new_n837_), .O(new_n917_));
  OR       g0901(.a(new_n917_), .b(new_n899_), .O(new_n918_));
  OR       g0902(.a(new_n918_), .b(new_n897_), .O(new_n919_));
  OR       g0903(.a(new_n919_), .b(new_n835_), .O(new_n920_));
  AND      g0904(.a(new_n920_), .b(i_2_6_62_0), .O(new_n921_));
  NOT      g0905(.a(new_n491_), .O(new_n922_));
  OR       g0906(.a(new_n482_), .b(new_n28_), .O(new_n923_));
  NAND     g0907(.a(new_n923_), .b(new_n278_), .O(new_n924_));
  AND      g0908(.a(new_n924_), .b(new_n605_), .O(new_n925_));
  AND      g0909(.a(new_n310_), .b(new_n230_), .O(new_n926_));
  OR       g0910(.a(new_n926_), .b(new_n925_), .O(new_n927_));
  AND      g0911(.a(new_n927_), .b(new_n456_), .O(new_n928_));
  AND      g0912(.a(new_n928_), .b(new_n922_), .O(new_n929_));
  OR       g0913(.a(new_n927_), .b(new_n193_), .O(new_n930_));
  AND      g0914(.a(new_n930_), .b(i_2_6_111_0), .O(new_n931_));
  AND      g0915(.a(new_n149_), .b(new_n193_), .O(new_n932_));
  OR       g0916(.a(new_n932_), .b(new_n928_), .O(new_n933_));
  AND      g0917(.a(new_n933_), .b(i_2_6_32_0), .O(new_n934_));
  OR       g0918(.a(new_n934_), .b(new_n931_), .O(new_n935_));
  AND      g0919(.a(new_n935_), .b(i_2_6_5_0), .O(new_n936_));
  OR       g0920(.a(new_n936_), .b(new_n929_), .O(new_n937_));
  AND      g0921(.a(new_n937_), .b(i_2_6_63_0), .O(new_n938_));
  OR       g0922(.a(new_n257_), .b(new_n23_), .O(new_n939_));
  AND      g0923(.a(new_n939_), .b(new_n68_), .O(new_n940_));
  AND      g0924(.a(new_n940_), .b(new_n747_), .O(new_n941_));
  OR       g0925(.a(new_n941_), .b(new_n938_), .O(new_n942_));
  AND      g0926(.a(new_n942_), .b(i_2_6_33_0), .O(new_n943_));
  OR       g0927(.a(new_n337_), .b(i_2_6_63_0), .O(new_n944_));
  AND      g0928(.a(new_n747_), .b(new_n114_), .O(new_n945_));
  AND      g0929(.a(new_n945_), .b(new_n944_), .O(new_n946_));
  OR       g0930(.a(new_n946_), .b(new_n943_), .O(new_n947_));
  AND      g0931(.a(new_n947_), .b(new_n35_), .O(new_n948_));
  OR       g0932(.a(new_n733_), .b(new_n324_), .O(new_n949_));
  AND      g0933(.a(new_n949_), .b(new_n23_), .O(new_n950_));
  AND      g0934(.a(new_n28_), .b(i_2_6_32_0), .O(new_n951_));
  AND      g0935(.a(new_n951_), .b(new_n278_), .O(new_n952_));
  OR       g0936(.a(new_n952_), .b(new_n338_), .O(new_n953_));
  AND      g0937(.a(new_n953_), .b(i_2_6_5_0), .O(new_n954_));
  OR       g0938(.a(new_n954_), .b(new_n385_), .O(new_n955_));
  OR       g0939(.a(new_n955_), .b(new_n950_), .O(new_n956_));
  AND      g0940(.a(new_n956_), .b(i_2_6_63_0), .O(new_n957_));
  AND      g0941(.a(new_n313_), .b(i_2_6_5_0), .O(new_n958_));
  AND      g0942(.a(new_n958_), .b(new_n339_), .O(new_n959_));
  OR       g0943(.a(new_n959_), .b(new_n957_), .O(new_n960_));
  AND      g0944(.a(new_n960_), .b(i_2_6_33_0), .O(new_n961_));
  OR       g0945(.a(new_n694_), .b(i_2_6_111_0), .O(new_n962_));
  AND      g0946(.a(new_n962_), .b(new_n19_), .O(new_n963_));
  OR       g0947(.a(new_n963_), .b(i_2_6_32_0), .O(new_n964_));
  AND      g0948(.a(new_n964_), .b(i_2_6_33_0), .O(new_n965_));
  AND      g0949(.a(new_n310_), .b(i_2_6_5_0), .O(new_n966_));
  NOT      g0950(.a(new_n527_), .O(new_n967_));
  NAND     g0951(.a(new_n967_), .b(new_n277_), .O(new_n968_));
  AND      g0952(.a(new_n968_), .b(new_n966_), .O(new_n969_));
  OR       g0953(.a(new_n969_), .b(new_n965_), .O(new_n970_));
  AND      g0954(.a(new_n970_), .b(i_2_6_63_0), .O(new_n971_));
  AND      g0955(.a(new_n733_), .b(new_n144_), .O(new_n972_));
  AND      g0956(.a(i_2_6_142_0), .b(i_2_6_120_0), .O(new_n973_));
  AND      g0957(.a(new_n973_), .b(i_2_6_110_0), .O(new_n974_));
  OR       g0958(.a(new_n974_), .b(new_n258_), .O(new_n975_));
  OR       g0959(.a(i_2_6_63_0), .b(i_2_6_5_0), .O(new_n976_));
  NOT      g0960(.a(new_n976_), .O(new_n977_));
  AND      g0961(.a(new_n977_), .b(new_n975_), .O(new_n978_));
  OR       g0962(.a(new_n978_), .b(new_n972_), .O(new_n979_));
  OR       g0963(.a(new_n584_), .b(new_n337_), .O(new_n980_));
  OR       g0964(.a(new_n980_), .b(new_n217_), .O(new_n981_));
  AND      g0965(.a(new_n981_), .b(i_2_6_33_0), .O(new_n982_));
  OR       g0966(.a(new_n319_), .b(i_2_6_33_0), .O(new_n983_));
  OR       g0967(.a(new_n983_), .b(new_n898_), .O(new_n984_));
  AND      g0968(.a(new_n984_), .b(i_2_6_5_0), .O(new_n985_));
  OR       g0969(.a(new_n985_), .b(new_n982_), .O(new_n986_));
  OR       g0970(.a(new_n986_), .b(new_n979_), .O(new_n987_));
  AND      g0971(.a(new_n987_), .b(new_n23_), .O(new_n988_));
  OR       g0972(.a(i_2_6_142_0), .b(i_2_6_111_0), .O(new_n989_));
  NAND     g0973(.a(new_n989_), .b(i_2_6_5_0), .O(new_n990_));
  OR       g0974(.a(new_n967_), .b(new_n276_), .O(new_n991_));
  NAND     g0975(.a(new_n991_), .b(new_n990_), .O(new_n992_));
  NAND     g0976(.a(new_n149_), .b(i_2_6_63_0), .O(new_n993_));
  OR       g0977(.a(i_2_6_124_0), .b(new_n463_), .O(new_n994_));
  OR       g0978(.a(new_n994_), .b(new_n736_), .O(new_n995_));
  NAND     g0979(.a(new_n995_), .b(new_n993_), .O(new_n996_));
  OR       g0980(.a(new_n996_), .b(new_n992_), .O(new_n997_));
  AND      g0981(.a(new_n997_), .b(i_2_6_32_0), .O(new_n998_));
  OR       g0982(.a(new_n998_), .b(new_n988_), .O(new_n999_));
  OR       g0983(.a(new_n999_), .b(new_n971_), .O(new_n1000_));
  AND      g0984(.a(new_n1000_), .b(new_n35_), .O(new_n1001_));
  AND      g0985(.a(new_n149_), .b(i_2_6_63_0), .O(new_n1002_));
  OR       g0986(.a(new_n1002_), .b(new_n127_), .O(new_n1003_));
  AND      g0987(.a(new_n34_), .b(i_2_6_5_0), .O(new_n1004_));
  AND      g0988(.a(new_n1004_), .b(new_n1003_), .O(new_n1005_));
  OR       g0989(.a(new_n1005_), .b(new_n1001_), .O(new_n1006_));
  OR       g0990(.a(new_n1006_), .b(new_n961_), .O(new_n1007_));
  AND      g0991(.a(new_n1007_), .b(new_n193_), .O(new_n1008_));
  NOT      g0992(.a(new_n310_), .O(new_n1009_));
  AND      g0993(.a(new_n1009_), .b(new_n217_), .O(new_n1010_));
  OR       g0994(.a(new_n1010_), .b(new_n46_), .O(new_n1011_));
  AND      g0995(.a(new_n1011_), .b(new_n722_), .O(new_n1012_));
  AND      g0996(.a(new_n645_), .b(i_2_6_63_0), .O(new_n1013_));
  OR       g0997(.a(new_n1013_), .b(new_n926_), .O(new_n1014_));
  AND      g0998(.a(new_n1014_), .b(new_n35_), .O(new_n1015_));
  AND      g0999(.a(new_n94_), .b(new_n694_), .O(new_n1016_));
  OR       g1000(.a(new_n1016_), .b(new_n217_), .O(new_n1017_));
  AND      g1001(.a(new_n1017_), .b(i_2_6_111_0), .O(new_n1018_));
  NAND     g1002(.a(new_n736_), .b(i_2_6_124_0), .O(new_n1019_));
  AND      g1003(.a(new_n1019_), .b(new_n78_), .O(new_n1020_));
  OR       g1004(.a(new_n1020_), .b(new_n1018_), .O(new_n1021_));
  OR       g1005(.a(new_n1021_), .b(new_n1015_), .O(new_n1022_));
  AND      g1006(.a(new_n1022_), .b(i_2_6_5_0), .O(new_n1023_));
  AND      g1007(.a(new_n394_), .b(i_2_6_63_0), .O(new_n1024_));
  AND      g1008(.a(new_n200_), .b(new_n109_), .O(new_n1025_));
  OR       g1009(.a(new_n1025_), .b(new_n1024_), .O(new_n1026_));
  OR       g1010(.a(new_n1026_), .b(new_n1023_), .O(new_n1027_));
  AND      g1011(.a(new_n1027_), .b(i_2_6_33_0), .O(new_n1028_));
  OR       g1012(.a(new_n1028_), .b(new_n1012_), .O(new_n1029_));
  AND      g1013(.a(new_n1029_), .b(i_2_6_32_0), .O(new_n1030_));
  AND      g1014(.a(new_n46_), .b(i_2_6_142_0), .O(new_n1031_));
  OR       g1015(.a(new_n1031_), .b(new_n966_), .O(new_n1032_));
  AND      g1016(.a(new_n1032_), .b(new_n95_), .O(new_n1033_));
  NOT      g1017(.a(new_n994_), .O(new_n1034_));
  AND      g1018(.a(new_n1034_), .b(new_n178_), .O(new_n1035_));
  OR       g1019(.a(new_n1035_), .b(new_n1033_), .O(new_n1036_));
  AND      g1020(.a(new_n1036_), .b(new_n557_), .O(new_n1037_));
  OR       g1021(.a(new_n1037_), .b(new_n1030_), .O(new_n1038_));
  OR       g1022(.a(new_n1038_), .b(new_n1008_), .O(new_n1039_));
  AND      g1023(.a(new_n1039_), .b(new_n18_), .O(new_n1040_));
  AND      g1024(.a(new_n217_), .b(i_2_6_33_0), .O(new_n1041_));
  AND      g1025(.a(new_n1041_), .b(new_n747_), .O(new_n1042_));
  AND      g1026(.a(new_n1042_), .b(new_n590_), .O(new_n1043_));
  OR       g1027(.a(new_n1043_), .b(new_n1040_), .O(new_n1044_));
  OR       g1028(.a(new_n1044_), .b(new_n948_), .O(new_n1045_));
  OR       g1029(.a(new_n1045_), .b(new_n921_), .O(new_n1046_));
  AND      g1030(.a(new_n1046_), .b(i_2_6_34_0), .O(new_n1047_));
  AND      g1031(.a(new_n338_), .b(new_n259_), .O(new_n1048_));
  NAND     g1032(.a(new_n923_), .b(new_n603_), .O(new_n1049_));
  OR       g1033(.a(new_n1049_), .b(new_n1048_), .O(new_n1050_));
  AND      g1034(.a(new_n1050_), .b(i_2_6_63_0), .O(new_n1051_));
  NOT      g1035(.a(new_n277_), .O(new_n1052_));
  AND      g1036(.a(new_n1052_), .b(new_n23_), .O(new_n1053_));
  OR       g1037(.a(new_n1053_), .b(new_n1051_), .O(new_n1054_));
  AND      g1038(.a(new_n1054_), .b(new_n18_), .O(new_n1055_));
  AND      g1039(.a(new_n206_), .b(new_n58_), .O(new_n1056_));
  OR       g1040(.a(new_n34_), .b(i_2_6_142_0), .O(new_n1057_));
  AND      g1041(.a(new_n1057_), .b(new_n199_), .O(new_n1058_));
  AND      g1042(.a(new_n354_), .b(i_2_6_111_0), .O(new_n1059_));
  OR       g1043(.a(new_n1059_), .b(new_n506_), .O(new_n1060_));
  AND      g1044(.a(new_n1060_), .b(new_n19_), .O(new_n1061_));
  OR       g1045(.a(new_n1061_), .b(new_n1058_), .O(new_n1062_));
  AND      g1046(.a(new_n1062_), .b(i_2_6_63_0), .O(new_n1063_));
  OR       g1047(.a(new_n1063_), .b(new_n1056_), .O(new_n1064_));
  AND      g1048(.a(new_n1064_), .b(i_2_6_62_0), .O(new_n1065_));
  OR       g1049(.a(new_n1065_), .b(new_n1055_), .O(new_n1066_));
  AND      g1050(.a(new_n1066_), .b(new_n193_), .O(new_n1067_));
  AND      g1051(.a(new_n313_), .b(new_n102_), .O(new_n1068_));
  NAND     g1052(.a(new_n775_), .b(new_n26_), .O(new_n1069_));
  AND      g1053(.a(new_n1069_), .b(new_n337_), .O(new_n1070_));
  AND      g1054(.a(new_n910_), .b(i_2_6_62_0), .O(new_n1071_));
  OR       g1055(.a(new_n1071_), .b(new_n1070_), .O(new_n1072_));
  AND      g1056(.a(new_n1072_), .b(i_2_6_142_0), .O(new_n1073_));
  OR       g1057(.a(new_n1073_), .b(new_n1068_), .O(new_n1074_));
  AND      g1058(.a(new_n1068_), .b(new_n140_), .O(new_n1075_));
  OR       g1059(.a(new_n1075_), .b(new_n23_), .O(new_n1076_));
  AND      g1060(.a(new_n1076_), .b(new_n452_), .O(new_n1077_));
  AND      g1061(.a(new_n1077_), .b(new_n1074_), .O(new_n1078_));
  OR       g1062(.a(new_n1078_), .b(new_n1067_), .O(new_n1079_));
  AND      g1063(.a(new_n1079_), .b(new_n35_), .O(new_n1080_));
  AND      g1064(.a(new_n337_), .b(i_2_6_32_0), .O(new_n1081_));
  OR       g1065(.a(new_n1081_), .b(new_n973_), .O(new_n1082_));
  NAND     g1066(.a(new_n1082_), .b(new_n95_), .O(new_n1083_));
  OR       g1067(.a(new_n923_), .b(new_n26_), .O(new_n1084_));
  NAND     g1068(.a(new_n1084_), .b(new_n1083_), .O(new_n1085_));
  AND      g1069(.a(new_n1085_), .b(i_2_6_111_0), .O(new_n1086_));
  NOT      g1070(.a(new_n236_), .O(new_n1087_));
  AND      g1071(.a(new_n491_), .b(new_n1087_), .O(new_n1088_));
  AND      g1072(.a(new_n1088_), .b(new_n195_), .O(new_n1089_));
  OR       g1073(.a(new_n1089_), .b(new_n1086_), .O(new_n1090_));
  AND      g1074(.a(new_n1090_), .b(new_n825_), .O(new_n1091_));
  OR       g1075(.a(new_n1091_), .b(new_n1080_), .O(new_n1092_));
  AND      g1076(.a(new_n1092_), .b(i_2_6_5_0), .O(new_n1093_));
  NOT      g1077(.a(new_n353_), .O(new_n1094_));
  OR       g1078(.a(new_n775_), .b(new_n26_), .O(new_n1095_));
  NAND     g1079(.a(new_n1095_), .b(new_n504_), .O(new_n1096_));
  AND      g1080(.a(new_n1096_), .b(new_n1094_), .O(new_n1097_));
  AND      g1081(.a(new_n582_), .b(new_n413_), .O(new_n1098_));
  OR       g1082(.a(new_n1098_), .b(new_n1097_), .O(new_n1099_));
  AND      g1083(.a(new_n1099_), .b(i_2_6_142_0), .O(new_n1100_));
  AND      g1084(.a(new_n932_), .b(new_n1052_), .O(new_n1101_));
  OR       g1085(.a(new_n1101_), .b(new_n1100_), .O(new_n1102_));
  AND      g1086(.a(new_n452_), .b(new_n41_), .O(new_n1103_));
  AND      g1087(.a(new_n1103_), .b(new_n1102_), .O(new_n1104_));
  OR       g1088(.a(new_n1104_), .b(new_n1093_), .O(new_n1105_));
  AND      g1089(.a(new_n1105_), .b(i_2_6_33_0), .O(new_n1106_));
  NOT      g1090(.a(new_n737_), .O(new_n1107_));
  AND      g1091(.a(new_n34_), .b(new_n366_), .O(new_n1108_));
  AND      g1092(.a(new_n1108_), .b(new_n1107_), .O(new_n1109_));
  AND      g1093(.a(new_n1109_), .b(new_n868_), .O(new_n1110_));
  OR       g1094(.a(new_n1110_), .b(new_n1106_), .O(new_n1111_));
  OR       g1095(.a(new_n1111_), .b(new_n1047_), .O(new_n1112_));
  OR       g1096(.a(new_n1112_), .b(new_n718_), .O(o_2_6_0_0));
endmodule


