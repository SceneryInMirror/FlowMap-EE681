// Benchmark "kernel_2_1" written by ABC on Wed May  4 16:37:49 2022

module kernel_2_1 ( 
    i_2_1_13_0, i_2_1_32_0, i_2_1_34_0, i_2_1_38_0, i_2_1_41_0, i_2_1_46_0,
    i_2_1_47_0, i_2_1_49_0, i_2_1_51_0, i_2_1_54_0, i_2_1_57_0, i_2_1_68_0,
    i_2_1_70_0, i_2_1_135_0, i_2_1_136_0,
    o_2_1_0_0  );
  input  i_2_1_13_0, i_2_1_32_0, i_2_1_34_0, i_2_1_38_0, i_2_1_41_0,
    i_2_1_46_0, i_2_1_47_0, i_2_1_49_0, i_2_1_51_0, i_2_1_54_0, i_2_1_57_0,
    i_2_1_68_0, i_2_1_70_0, i_2_1_135_0, i_2_1_136_0;
  output o_2_1_0_0;
  wire new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_, new_n1329_, new_n1330_,
    new_n1331_, new_n1332_, new_n1333_, new_n1334_, new_n1335_, new_n1336_,
    new_n1337_, new_n1338_, new_n1339_, new_n1340_, new_n1341_, new_n1342_,
    new_n1343_, new_n1344_, new_n1345_, new_n1346_, new_n1347_, new_n1348_,
    new_n1349_, new_n1350_, new_n1351_, new_n1352_, new_n1353_, new_n1354_,
    new_n1355_, new_n1356_, new_n1357_, new_n1358_, new_n1359_, new_n1360_,
    new_n1361_, new_n1362_, new_n1363_, new_n1364_, new_n1365_, new_n1366_,
    new_n1367_, new_n1368_, new_n1369_, new_n1370_, new_n1371_, new_n1372_,
    new_n1373_, new_n1374_, new_n1375_, new_n1376_, new_n1377_, new_n1378_,
    new_n1379_, new_n1380_, new_n1381_, new_n1382_, new_n1383_, new_n1384_,
    new_n1385_, new_n1386_, new_n1387_, new_n1388_, new_n1389_, new_n1390_,
    new_n1391_, new_n1392_, new_n1393_, new_n1394_, new_n1395_, new_n1396_,
    new_n1397_, new_n1398_, new_n1399_, new_n1400_, new_n1401_, new_n1402_,
    new_n1403_, new_n1404_, new_n1405_, new_n1406_, new_n1407_, new_n1408_,
    new_n1409_, new_n1410_, new_n1411_, new_n1412_, new_n1413_, new_n1414_,
    new_n1415_, new_n1416_, new_n1417_, new_n1418_, new_n1419_, new_n1420_,
    new_n1421_, new_n1422_, new_n1423_, new_n1424_, new_n1425_, new_n1426_,
    new_n1427_, new_n1428_, new_n1429_, new_n1430_, new_n1431_, new_n1432_,
    new_n1433_, new_n1434_, new_n1435_, new_n1436_, new_n1437_, new_n1438_,
    new_n1439_, new_n1440_, new_n1441_, new_n1442_, new_n1443_, new_n1444_,
    new_n1445_, new_n1446_, new_n1447_, new_n1448_, new_n1449_, new_n1450_,
    new_n1451_, new_n1452_, new_n1453_, new_n1454_, new_n1455_, new_n1456_,
    new_n1457_, new_n1458_, new_n1459_, new_n1460_, new_n1461_, new_n1462_,
    new_n1463_, new_n1464_, new_n1465_, new_n1466_, new_n1467_, new_n1468_,
    new_n1469_, new_n1470_, new_n1471_, new_n1472_, new_n1473_, new_n1474_,
    new_n1475_, new_n1476_, new_n1477_, new_n1478_, new_n1479_, new_n1480_,
    new_n1481_, new_n1482_, new_n1483_, new_n1484_, new_n1485_, new_n1486_,
    new_n1487_, new_n1488_, new_n1489_, new_n1490_, new_n1491_, new_n1492_,
    new_n1493_, new_n1494_, new_n1495_, new_n1496_, new_n1497_, new_n1498_,
    new_n1499_, new_n1500_, new_n1501_, new_n1502_, new_n1503_, new_n1504_,
    new_n1505_, new_n1506_, new_n1507_, new_n1508_, new_n1509_, new_n1510_,
    new_n1511_, new_n1512_, new_n1513_, new_n1514_, new_n1515_, new_n1516_,
    new_n1517_, new_n1518_, new_n1519_, new_n1520_, new_n1521_, new_n1522_,
    new_n1523_, new_n1524_, new_n1525_, new_n1526_, new_n1527_, new_n1528_,
    new_n1529_, new_n1530_, new_n1531_, new_n1532_, new_n1533_, new_n1534_,
    new_n1535_, new_n1536_, new_n1537_, new_n1538_, new_n1539_, new_n1540_,
    new_n1541_, new_n1542_, new_n1543_, new_n1544_, new_n1545_, new_n1546_,
    new_n1547_, new_n1548_, new_n1549_, new_n1550_, new_n1551_, new_n1552_,
    new_n1553_, new_n1554_, new_n1555_, new_n1556_, new_n1557_, new_n1558_,
    new_n1559_, new_n1560_, new_n1561_, new_n1562_, new_n1563_, new_n1564_,
    new_n1565_, new_n1566_, new_n1567_, new_n1568_, new_n1569_, new_n1570_,
    new_n1571_, new_n1572_, new_n1573_, new_n1574_, new_n1575_, new_n1576_,
    new_n1577_, new_n1578_, new_n1579_, new_n1580_, new_n1581_, new_n1582_,
    new_n1583_, new_n1584_, new_n1585_, new_n1586_, new_n1587_, new_n1588_,
    new_n1589_, new_n1590_, new_n1591_, new_n1592_, new_n1593_, new_n1594_,
    new_n1595_, new_n1596_, new_n1597_, new_n1598_, new_n1599_, new_n1600_,
    new_n1601_, new_n1602_, new_n1603_, new_n1604_, new_n1605_, new_n1606_,
    new_n1607_, new_n1608_, new_n1609_, new_n1610_, new_n1611_, new_n1612_,
    new_n1613_, new_n1614_, new_n1615_, new_n1616_, new_n1617_, new_n1618_,
    new_n1619_, new_n1620_, new_n1621_, new_n1622_, new_n1623_, new_n1624_,
    new_n1625_, new_n1626_, new_n1627_, new_n1628_, new_n1629_, new_n1630_,
    new_n1631_, new_n1632_, new_n1633_, new_n1634_, new_n1635_, new_n1636_,
    new_n1637_, new_n1638_, new_n1639_, new_n1640_, new_n1641_, new_n1642_,
    new_n1643_, new_n1644_, new_n1645_, new_n1646_, new_n1647_, new_n1648_,
    new_n1649_, new_n1650_, new_n1651_, new_n1652_, new_n1653_, new_n1654_,
    new_n1655_, new_n1656_, new_n1657_, new_n1658_, new_n1659_, new_n1660_,
    new_n1661_, new_n1662_, new_n1663_, new_n1664_, new_n1665_, new_n1666_,
    new_n1667_, new_n1668_, new_n1669_, new_n1670_, new_n1671_, new_n1672_,
    new_n1673_, new_n1674_, new_n1675_, new_n1676_, new_n1677_, new_n1678_,
    new_n1679_, new_n1680_, new_n1681_, new_n1682_, new_n1683_, new_n1684_,
    new_n1685_, new_n1686_, new_n1687_, new_n1688_, new_n1689_, new_n1690_,
    new_n1691_, new_n1692_, new_n1693_, new_n1694_, new_n1695_, new_n1696_,
    new_n1697_, new_n1698_, new_n1699_, new_n1700_, new_n1701_, new_n1702_,
    new_n1703_, new_n1704_, new_n1705_, new_n1706_, new_n1707_, new_n1708_,
    new_n1709_, new_n1710_, new_n1711_, new_n1712_, new_n1713_, new_n1714_,
    new_n1715_, new_n1716_, new_n1717_, new_n1718_, new_n1719_, new_n1720_,
    new_n1721_, new_n1722_, new_n1723_, new_n1724_, new_n1725_, new_n1726_,
    new_n1727_, new_n1728_, new_n1729_, new_n1730_, new_n1731_, new_n1732_,
    new_n1733_, new_n1734_, new_n1735_, new_n1736_, new_n1737_, new_n1738_,
    new_n1739_, new_n1740_, new_n1741_, new_n1742_, new_n1743_, new_n1744_,
    new_n1745_, new_n1746_, new_n1747_, new_n1748_, new_n1749_, new_n1750_,
    new_n1751_, new_n1752_, new_n1753_, new_n1754_, new_n1755_, new_n1756_,
    new_n1757_, new_n1758_, new_n1759_, new_n1760_, new_n1761_, new_n1762_,
    new_n1763_, new_n1764_, new_n1765_, new_n1766_, new_n1767_, new_n1768_,
    new_n1769_, new_n1770_, new_n1771_, new_n1772_, new_n1773_, new_n1774_,
    new_n1775_, new_n1776_, new_n1777_, new_n1778_, new_n1779_, new_n1780_,
    new_n1781_, new_n1782_, new_n1783_, new_n1784_, new_n1785_, new_n1786_,
    new_n1787_, new_n1788_, new_n1789_, new_n1790_, new_n1791_, new_n1792_,
    new_n1793_, new_n1794_, new_n1795_, new_n1796_, new_n1797_, new_n1798_,
    new_n1799_, new_n1800_, new_n1801_, new_n1802_, new_n1803_, new_n1804_,
    new_n1805_, new_n1806_, new_n1807_, new_n1808_, new_n1809_, new_n1810_,
    new_n1811_, new_n1812_, new_n1813_, new_n1814_, new_n1815_, new_n1816_,
    new_n1817_, new_n1818_, new_n1819_, new_n1820_, new_n1821_, new_n1822_,
    new_n1823_, new_n1824_, new_n1825_, new_n1826_, new_n1827_, new_n1828_,
    new_n1829_, new_n1830_, new_n1831_, new_n1832_, new_n1833_, new_n1834_,
    new_n1835_, new_n1836_, new_n1837_, new_n1838_, new_n1839_, new_n1840_,
    new_n1841_, new_n1842_, new_n1843_, new_n1844_, new_n1845_, new_n1846_,
    new_n1847_, new_n1848_, new_n1849_, new_n1850_, new_n1851_, new_n1852_,
    new_n1853_, new_n1854_, new_n1855_, new_n1856_, new_n1857_, new_n1858_,
    new_n1859_, new_n1860_, new_n1861_, new_n1862_, new_n1863_, new_n1864_,
    new_n1865_, new_n1866_, new_n1867_, new_n1868_, new_n1869_, new_n1870_,
    new_n1871_, new_n1872_, new_n1873_, new_n1874_, new_n1875_, new_n1876_,
    new_n1877_, new_n1878_, new_n1879_, new_n1880_, new_n1881_, new_n1882_,
    new_n1883_, new_n1884_, new_n1885_, new_n1886_, new_n1887_, new_n1888_,
    new_n1889_, new_n1890_, new_n1891_, new_n1892_, new_n1893_, new_n1894_,
    new_n1895_, new_n1896_, new_n1897_, new_n1898_, new_n1899_, new_n1900_,
    new_n1901_, new_n1902_, new_n1903_, new_n1904_, new_n1905_, new_n1906_,
    new_n1907_, new_n1908_, new_n1909_, new_n1910_, new_n1911_, new_n1912_,
    new_n1913_, new_n1914_, new_n1915_, new_n1916_, new_n1917_, new_n1918_,
    new_n1919_, new_n1920_, new_n1921_, new_n1922_, new_n1923_, new_n1924_,
    new_n1925_, new_n1926_, new_n1927_, new_n1928_, new_n1929_, new_n1930_,
    new_n1931_, new_n1932_, new_n1933_, new_n1934_, new_n1935_, new_n1936_,
    new_n1937_, new_n1938_, new_n1939_, new_n1940_, new_n1941_, new_n1942_,
    new_n1943_, new_n1944_, new_n1945_, new_n1946_, new_n1947_, new_n1948_,
    new_n1949_, new_n1950_, new_n1951_, new_n1952_, new_n1953_, new_n1954_,
    new_n1955_, new_n1956_, new_n1957_, new_n1958_, new_n1959_, new_n1960_,
    new_n1961_, new_n1962_, new_n1963_, new_n1964_, new_n1965_, new_n1966_,
    new_n1967_, new_n1968_, new_n1969_, new_n1970_, new_n1971_, new_n1972_,
    new_n1973_, new_n1974_, new_n1975_, new_n1976_, new_n1977_, new_n1978_,
    new_n1979_, new_n1980_, new_n1981_, new_n1982_, new_n1983_, new_n1984_,
    new_n1985_, new_n1986_, new_n1987_, new_n1988_, new_n1989_, new_n1990_,
    new_n1991_, new_n1992_, new_n1993_, new_n1994_, new_n1995_, new_n1996_,
    new_n1997_, new_n1998_, new_n1999_, new_n2000_, new_n2001_, new_n2002_,
    new_n2003_, new_n2004_, new_n2005_, new_n2006_, new_n2007_, new_n2008_,
    new_n2009_, new_n2010_, new_n2011_, new_n2012_, new_n2013_, new_n2014_,
    new_n2015_, new_n2016_, new_n2017_, new_n2018_, new_n2019_, new_n2020_,
    new_n2021_, new_n2022_, new_n2023_, new_n2024_, new_n2025_, new_n2026_,
    new_n2027_, new_n2028_, new_n2029_, new_n2030_, new_n2031_, new_n2032_,
    new_n2033_, new_n2034_, new_n2035_, new_n2036_, new_n2037_, new_n2038_,
    new_n2039_, new_n2040_, new_n2041_, new_n2042_, new_n2043_, new_n2044_,
    new_n2045_, new_n2046_, new_n2047_, new_n2048_, new_n2049_, new_n2050_,
    new_n2051_, new_n2052_, new_n2053_, new_n2054_, new_n2055_, new_n2056_,
    new_n2057_, new_n2058_, new_n2059_, new_n2060_, new_n2061_, new_n2062_,
    new_n2063_, new_n2064_, new_n2065_, new_n2066_, new_n2067_, new_n2068_,
    new_n2069_, new_n2070_, new_n2071_, new_n2072_, new_n2073_, new_n2074_,
    new_n2075_, new_n2076_, new_n2077_, new_n2078_, new_n2079_, new_n2080_,
    new_n2081_, new_n2082_, new_n2083_, new_n2084_, new_n2085_, new_n2086_,
    new_n2087_, new_n2088_, new_n2089_, new_n2090_, new_n2091_, new_n2092_,
    new_n2093_, new_n2094_, new_n2095_, new_n2096_, new_n2097_, new_n2098_,
    new_n2099_, new_n2100_, new_n2101_, new_n2102_, new_n2103_, new_n2104_,
    new_n2105_, new_n2106_, new_n2107_, new_n2108_, new_n2109_, new_n2110_,
    new_n2111_, new_n2112_, new_n2113_, new_n2114_, new_n2115_, new_n2116_,
    new_n2117_, new_n2118_, new_n2119_, new_n2120_, new_n2121_, new_n2122_,
    new_n2123_, new_n2124_, new_n2125_, new_n2126_, new_n2127_, new_n2128_,
    new_n2129_, new_n2130_, new_n2131_, new_n2132_, new_n2133_, new_n2134_,
    new_n2135_, new_n2136_, new_n2137_, new_n2138_, new_n2139_, new_n2140_,
    new_n2141_, new_n2142_, new_n2143_, new_n2144_, new_n2145_, new_n2146_,
    new_n2147_, new_n2148_, new_n2149_, new_n2150_, new_n2151_, new_n2152_,
    new_n2153_, new_n2154_, new_n2155_, new_n2156_, new_n2157_, new_n2158_,
    new_n2159_, new_n2160_, new_n2161_, new_n2162_, new_n2163_, new_n2164_,
    new_n2165_, new_n2166_, new_n2167_, new_n2168_, new_n2169_, new_n2170_,
    new_n2171_, new_n2172_, new_n2173_, new_n2174_, new_n2175_, new_n2176_,
    new_n2177_, new_n2178_, new_n2179_, new_n2180_, new_n2181_, new_n2182_,
    new_n2183_, new_n2184_, new_n2185_, new_n2186_, new_n2187_, new_n2188_,
    new_n2189_, new_n2190_, new_n2191_, new_n2192_, new_n2193_, new_n2194_,
    new_n2195_, new_n2196_, new_n2197_, new_n2198_, new_n2199_, new_n2200_,
    new_n2201_, new_n2202_, new_n2203_, new_n2204_, new_n2205_, new_n2206_,
    new_n2207_, new_n2208_, new_n2209_, new_n2210_, new_n2211_, new_n2212_,
    new_n2213_, new_n2214_, new_n2215_, new_n2216_, new_n2217_, new_n2218_,
    new_n2219_, new_n2220_, new_n2221_, new_n2222_, new_n2223_, new_n2224_,
    new_n2225_;
  NOT      g0000(.a(i_2_1_47_0), .O(new_n17_));
  NOT      g0001(.a(i_2_1_51_0), .O(new_n18_));
  NOT      g0002(.a(i_2_1_46_0), .O(new_n19_));
  NOT      g0003(.a(i_2_1_57_0), .O(new_n20_));
  AND      g0004(.a(i_2_1_136_0), .b(i_2_1_135_0), .O(new_n21_));
  OR       g0005(.a(new_n21_), .b(i_2_1_70_0), .O(new_n22_));
  AND      g0006(.a(new_n22_), .b(i_2_1_68_0), .O(new_n23_));
  OR       g0007(.a(new_n23_), .b(new_n20_), .O(new_n24_));
  NOT      g0008(.a(i_2_1_68_0), .O(new_n25_));
  OR       g0009(.a(new_n25_), .b(i_2_1_49_0), .O(new_n26_));
  NOT      g0010(.a(i_2_1_136_0), .O(new_n27_));
  OR       g0011(.a(new_n27_), .b(i_2_1_49_0), .O(new_n28_));
  OR       g0012(.a(new_n28_), .b(i_2_1_135_0), .O(new_n29_));
  NAND     g0013(.a(new_n29_), .b(new_n26_), .O(new_n30_));
  AND      g0014(.a(new_n30_), .b(new_n24_), .O(new_n31_));
  NOT      g0015(.a(i_2_1_54_0), .O(new_n32_));
  OR       g0016(.a(i_2_1_70_0), .b(i_2_1_49_0), .O(new_n33_));
  NAND     g0017(.a(i_2_1_70_0), .b(i_2_1_34_0), .O(new_n34_));
  NAND     g0018(.a(new_n34_), .b(new_n33_), .O(new_n35_));
  AND      g0019(.a(new_n35_), .b(new_n32_), .O(new_n36_));
  AND      g0020(.a(i_2_1_70_0), .b(i_2_1_68_0), .O(new_n37_));
  AND      g0021(.a(new_n37_), .b(i_2_1_136_0), .O(new_n38_));
  AND      g0022(.a(i_2_1_136_0), .b(i_2_1_68_0), .O(new_n39_));
  OR       g0023(.a(new_n39_), .b(new_n20_), .O(new_n40_));
  AND      g0024(.a(new_n40_), .b(i_2_1_13_0), .O(new_n41_));
  OR       g0025(.a(new_n41_), .b(new_n38_), .O(new_n42_));
  OR       g0026(.a(new_n42_), .b(new_n36_), .O(new_n43_));
  OR       g0027(.a(i_2_1_70_0), .b(i_2_1_68_0), .O(new_n44_));
  AND      g0028(.a(new_n44_), .b(i_2_1_135_0), .O(new_n45_));
  OR       g0029(.a(new_n27_), .b(i_2_1_57_0), .O(new_n46_));
  OR       g0030(.a(i_2_1_68_0), .b(i_2_1_38_0), .O(new_n47_));
  NAND     g0031(.a(new_n47_), .b(i_2_1_70_0), .O(new_n48_));
  NAND     g0032(.a(new_n48_), .b(new_n46_), .O(new_n49_));
  NAND     g0033(.a(new_n49_), .b(new_n45_), .O(new_n50_));
  AND      g0034(.a(i_2_1_70_0), .b(i_2_1_49_0), .O(new_n51_));
  NOT      g0035(.a(i_2_1_34_0), .O(new_n52_));
  NOT      g0036(.a(i_2_1_70_0), .O(new_n53_));
  NOT      g0037(.a(i_2_1_135_0), .O(new_n54_));
  OR       g0038(.a(i_2_1_136_0), .b(new_n54_), .O(new_n55_));
  AND      g0039(.a(new_n55_), .b(new_n53_), .O(new_n56_));
  OR       g0040(.a(new_n56_), .b(new_n52_), .O(new_n57_));
  OR       g0041(.a(new_n57_), .b(new_n51_), .O(new_n58_));
  NAND     g0042(.a(new_n58_), .b(new_n50_), .O(new_n59_));
  OR       g0043(.a(new_n59_), .b(new_n43_), .O(new_n60_));
  OR       g0044(.a(new_n60_), .b(new_n31_), .O(new_n61_));
  AND      g0045(.a(new_n61_), .b(i_2_1_41_0), .O(new_n62_));
  NOT      g0046(.a(i_2_1_49_0), .O(new_n63_));
  AND      g0047(.a(new_n32_), .b(i_2_1_34_0), .O(new_n64_));
  OR       g0048(.a(i_2_1_135_0), .b(new_n20_), .O(new_n65_));
  OR       g0049(.a(new_n65_), .b(i_2_1_136_0), .O(new_n66_));
  OR       g0050(.a(new_n66_), .b(new_n64_), .O(new_n67_));
  OR       g0051(.a(i_2_1_70_0), .b(i_2_1_38_0), .O(new_n68_));
  OR       g0052(.a(new_n64_), .b(i_2_1_68_0), .O(new_n69_));
  AND      g0053(.a(new_n69_), .b(new_n68_), .O(new_n70_));
  AND      g0054(.a(new_n70_), .b(new_n67_), .O(new_n71_));
  OR       g0055(.a(i_2_1_68_0), .b(new_n32_), .O(new_n72_));
  AND      g0056(.a(i_2_1_70_0), .b(i_2_1_38_0), .O(new_n73_));
  AND      g0057(.a(i_2_1_135_0), .b(i_2_1_34_0), .O(new_n74_));
  OR       g0058(.a(new_n74_), .b(new_n73_), .O(new_n75_));
  AND      g0059(.a(new_n75_), .b(new_n72_), .O(new_n76_));
  AND      g0060(.a(i_2_1_68_0), .b(new_n20_), .O(new_n77_));
  AND      g0061(.a(new_n77_), .b(new_n21_), .O(new_n78_));
  OR       g0062(.a(i_2_1_57_0), .b(i_2_1_54_0), .O(new_n79_));
  NOT      g0063(.a(new_n79_), .O(new_n80_));
  OR       g0064(.a(new_n80_), .b(new_n78_), .O(new_n81_));
  AND      g0065(.a(i_2_1_135_0), .b(i_2_1_38_0), .O(new_n82_));
  NAND     g0066(.a(new_n82_), .b(i_2_1_136_0), .O(new_n83_));
  OR       g0067(.a(i_2_1_135_0), .b(i_2_1_70_0), .O(new_n84_));
  NOT      g0068(.a(new_n84_), .O(new_n85_));
  OR       g0069(.a(new_n25_), .b(i_2_1_54_0), .O(new_n86_));
  OR       g0070(.a(new_n86_), .b(new_n85_), .O(new_n87_));
  NAND     g0071(.a(new_n87_), .b(new_n83_), .O(new_n88_));
  OR       g0072(.a(new_n88_), .b(new_n81_), .O(new_n89_));
  OR       g0073(.a(new_n89_), .b(new_n76_), .O(new_n90_));
  OR       g0074(.a(new_n90_), .b(new_n71_), .O(new_n91_));
  AND      g0075(.a(new_n91_), .b(new_n63_), .O(new_n92_));
  OR       g0076(.a(i_2_1_70_0), .b(new_n20_), .O(new_n93_));
  OR       g0077(.a(i_2_1_135_0), .b(new_n63_), .O(new_n94_));
  AND      g0078(.a(new_n94_), .b(new_n93_), .O(new_n95_));
  OR       g0079(.a(i_2_1_136_0), .b(new_n63_), .O(new_n96_));
  AND      g0080(.a(new_n96_), .b(i_2_1_135_0), .O(new_n97_));
  NAND     g0081(.a(new_n46_), .b(i_2_1_54_0), .O(new_n98_));
  OR       g0082(.a(new_n98_), .b(new_n97_), .O(new_n99_));
  OR       g0083(.a(new_n99_), .b(new_n95_), .O(new_n100_));
  AND      g0084(.a(new_n100_), .b(i_2_1_68_0), .O(new_n101_));
  NOT      g0085(.a(i_2_1_38_0), .O(new_n102_));
  AND      g0086(.a(i_2_1_135_0), .b(i_2_1_68_0), .O(new_n103_));
  NOT      g0087(.a(new_n103_), .O(new_n104_));
  AND      g0088(.a(new_n104_), .b(i_2_1_49_0), .O(new_n105_));
  OR       g0089(.a(new_n105_), .b(new_n102_), .O(new_n106_));
  NAND     g0090(.a(new_n72_), .b(i_2_1_34_0), .O(new_n107_));
  NAND     g0091(.a(new_n107_), .b(new_n106_), .O(new_n108_));
  OR       g0092(.a(new_n108_), .b(new_n101_), .O(new_n109_));
  AND      g0093(.a(new_n109_), .b(i_2_1_13_0), .O(new_n110_));
  OR       g0094(.a(new_n54_), .b(i_2_1_54_0), .O(new_n111_));
  OR       g0095(.a(new_n111_), .b(new_n53_), .O(new_n112_));
  OR       g0096(.a(new_n27_), .b(i_2_1_54_0), .O(new_n113_));
  OR       g0097(.a(new_n113_), .b(new_n54_), .O(new_n114_));
  AND      g0098(.a(new_n114_), .b(new_n86_), .O(new_n115_));
  NAND     g0099(.a(new_n115_), .b(new_n112_), .O(new_n116_));
  NAND     g0100(.a(new_n22_), .b(i_2_1_68_0), .O(new_n117_));
  AND      g0101(.a(new_n111_), .b(new_n27_), .O(new_n118_));
  OR       g0102(.a(new_n118_), .b(i_2_1_57_0), .O(new_n119_));
  NAND     g0103(.a(new_n119_), .b(new_n117_), .O(new_n120_));
  OR       g0104(.a(new_n120_), .b(new_n116_), .O(new_n121_));
  AND      g0105(.a(new_n121_), .b(i_2_1_34_0), .O(new_n122_));
  AND      g0106(.a(i_2_1_135_0), .b(i_2_1_70_0), .O(new_n123_));
  AND      g0107(.a(new_n123_), .b(i_2_1_136_0), .O(new_n124_));
  AND      g0108(.a(new_n20_), .b(i_2_1_38_0), .O(new_n125_));
  AND      g0109(.a(new_n125_), .b(new_n124_), .O(new_n126_));
  OR       g0110(.a(i_2_1_136_0), .b(i_2_1_135_0), .O(new_n127_));
  AND      g0111(.a(i_2_1_70_0), .b(new_n20_), .O(new_n128_));
  AND      g0112(.a(new_n128_), .b(new_n127_), .O(new_n129_));
  OR       g0113(.a(new_n129_), .b(new_n32_), .O(new_n130_));
  AND      g0114(.a(new_n103_), .b(i_2_1_136_0), .O(new_n131_));
  OR       g0115(.a(new_n131_), .b(new_n77_), .O(new_n132_));
  AND      g0116(.a(new_n132_), .b(new_n130_), .O(new_n133_));
  OR       g0117(.a(new_n133_), .b(new_n126_), .O(new_n134_));
  OR       g0118(.a(new_n134_), .b(new_n122_), .O(new_n135_));
  OR       g0119(.a(new_n135_), .b(new_n110_), .O(new_n136_));
  OR       g0120(.a(new_n136_), .b(new_n92_), .O(new_n137_));
  OR       g0121(.a(new_n137_), .b(new_n62_), .O(new_n138_));
  AND      g0122(.a(new_n138_), .b(new_n19_), .O(new_n139_));
  OR       g0123(.a(new_n32_), .b(i_2_1_13_0), .O(new_n140_));
  AND      g0124(.a(new_n63_), .b(i_2_1_34_0), .O(new_n141_));
  OR       g0125(.a(new_n141_), .b(new_n68_), .O(new_n142_));
  OR       g0126(.a(new_n142_), .b(new_n140_), .O(new_n143_));
  AND      g0127(.a(new_n69_), .b(new_n63_), .O(new_n144_));
  NAND     g0128(.a(new_n144_), .b(new_n143_), .O(new_n145_));
  NAND     g0129(.a(new_n145_), .b(new_n34_), .O(new_n146_));
  AND      g0130(.a(new_n146_), .b(i_2_1_136_0), .O(new_n147_));
  AND      g0131(.a(i_2_1_136_0), .b(new_n63_), .O(new_n148_));
  OR       g0132(.a(new_n148_), .b(i_2_1_70_0), .O(new_n149_));
  OR       g0133(.a(new_n149_), .b(new_n32_), .O(new_n150_));
  AND      g0134(.a(new_n150_), .b(new_n69_), .O(new_n151_));
  OR       g0135(.a(new_n27_), .b(i_2_1_68_0), .O(new_n152_));
  AND      g0136(.a(new_n96_), .b(i_2_1_13_0), .O(new_n153_));
  AND      g0137(.a(new_n153_), .b(new_n152_), .O(new_n154_));
  OR       g0138(.a(new_n19_), .b(i_2_1_34_0), .O(new_n155_));
  OR       g0139(.a(new_n155_), .b(i_2_1_136_0), .O(new_n156_));
  NAND     g0140(.a(new_n156_), .b(i_2_1_54_0), .O(new_n157_));
  AND      g0141(.a(new_n157_), .b(i_2_1_38_0), .O(new_n158_));
  OR       g0142(.a(new_n158_), .b(new_n154_), .O(new_n159_));
  OR       g0143(.a(new_n159_), .b(new_n151_), .O(new_n160_));
  AND      g0144(.a(new_n160_), .b(new_n20_), .O(new_n161_));
  OR       g0145(.a(new_n161_), .b(new_n147_), .O(new_n162_));
  AND      g0146(.a(new_n162_), .b(i_2_1_135_0), .O(new_n163_));
  OR       g0147(.a(new_n27_), .b(i_2_1_135_0), .O(new_n164_));
  NAND     g0148(.a(new_n164_), .b(new_n53_), .O(new_n165_));
  AND      g0149(.a(new_n165_), .b(new_n31_), .O(new_n166_));
  OR       g0150(.a(new_n32_), .b(i_2_1_34_0), .O(new_n167_));
  NAND     g0151(.a(new_n167_), .b(i_2_1_68_0), .O(new_n168_));
  AND      g0152(.a(i_2_1_57_0), .b(i_2_1_49_0), .O(new_n169_));
  OR       g0153(.a(new_n169_), .b(new_n102_), .O(new_n170_));
  NAND     g0154(.a(new_n170_), .b(new_n168_), .O(new_n171_));
  OR       g0155(.a(new_n171_), .b(new_n166_), .O(new_n172_));
  AND      g0156(.a(new_n172_), .b(i_2_1_13_0), .O(new_n173_));
  NAND     g0157(.a(new_n77_), .b(i_2_1_70_0), .O(new_n174_));
  AND      g0158(.a(new_n27_), .b(i_2_1_135_0), .O(new_n175_));
  AND      g0159(.a(i_2_1_68_0), .b(i_2_1_13_0), .O(new_n176_));
  AND      g0160(.a(new_n176_), .b(new_n175_), .O(new_n177_));
  AND      g0161(.a(i_2_1_136_0), .b(new_n32_), .O(new_n178_));
  AND      g0162(.a(new_n178_), .b(new_n54_), .O(new_n179_));
  OR       g0163(.a(new_n179_), .b(new_n177_), .O(new_n180_));
  NAND     g0164(.a(new_n180_), .b(i_2_1_57_0), .O(new_n181_));
  NAND     g0165(.a(new_n181_), .b(new_n174_), .O(new_n182_));
  AND      g0166(.a(new_n182_), .b(i_2_1_49_0), .O(new_n183_));
  AND      g0167(.a(new_n98_), .b(i_2_1_68_0), .O(new_n184_));
  AND      g0168(.a(new_n141_), .b(new_n72_), .O(new_n185_));
  OR       g0169(.a(new_n185_), .b(new_n178_), .O(new_n186_));
  OR       g0170(.a(new_n186_), .b(new_n184_), .O(new_n187_));
  AND      g0171(.a(new_n187_), .b(i_2_1_70_0), .O(new_n188_));
  OR       g0172(.a(i_2_1_57_0), .b(i_2_1_49_0), .O(new_n189_));
  NOT      g0173(.a(new_n189_), .O(new_n190_));
  AND      g0174(.a(new_n190_), .b(i_2_1_68_0), .O(new_n191_));
  AND      g0175(.a(i_2_1_68_0), .b(new_n63_), .O(new_n192_));
  OR       g0176(.a(i_2_1_136_0), .b(i_2_1_57_0), .O(new_n193_));
  NOT      g0177(.a(new_n193_), .O(new_n194_));
  OR       g0178(.a(new_n194_), .b(new_n192_), .O(new_n195_));
  AND      g0179(.a(new_n195_), .b(i_2_1_34_0), .O(new_n196_));
  OR       g0180(.a(new_n196_), .b(new_n191_), .O(new_n197_));
  AND      g0181(.a(new_n197_), .b(new_n32_), .O(new_n198_));
  NOT      g0182(.a(new_n46_), .O(new_n199_));
  AND      g0183(.a(new_n199_), .b(i_2_1_68_0), .O(new_n200_));
  OR       g0184(.a(new_n200_), .b(new_n141_), .O(new_n201_));
  AND      g0185(.a(new_n201_), .b(i_2_1_38_0), .O(new_n202_));
  OR       g0186(.a(new_n202_), .b(new_n198_), .O(new_n203_));
  OR       g0187(.a(new_n203_), .b(new_n188_), .O(new_n204_));
  OR       g0188(.a(new_n204_), .b(new_n183_), .O(new_n205_));
  OR       g0189(.a(new_n205_), .b(new_n173_), .O(new_n206_));
  OR       g0190(.a(new_n206_), .b(new_n163_), .O(new_n207_));
  AND      g0191(.a(new_n207_), .b(i_2_1_41_0), .O(new_n208_));
  OR       g0192(.a(i_2_1_135_0), .b(i_2_1_68_0), .O(new_n209_));
  NAND     g0193(.a(new_n209_), .b(new_n105_), .O(new_n210_));
  AND      g0194(.a(new_n210_), .b(i_2_1_13_0), .O(new_n211_));
  AND      g0195(.a(i_2_1_136_0), .b(i_2_1_34_0), .O(new_n212_));
  OR       g0196(.a(new_n212_), .b(new_n192_), .O(new_n213_));
  AND      g0197(.a(new_n213_), .b(new_n32_), .O(new_n214_));
  AND      g0198(.a(new_n54_), .b(i_2_1_68_0), .O(new_n215_));
  OR       g0199(.a(new_n215_), .b(i_2_1_34_0), .O(new_n216_));
  AND      g0200(.a(new_n216_), .b(i_2_1_70_0), .O(new_n217_));
  NAND     g0201(.a(i_2_1_136_0), .b(i_2_1_135_0), .O(new_n218_));
  OR       g0202(.a(new_n26_), .b(new_n218_), .O(new_n219_));
  NOT      g0203(.a(i_2_1_41_0), .O(new_n220_));
  NAND     g0204(.a(new_n74_), .b(new_n220_), .O(new_n221_));
  NAND     g0205(.a(new_n221_), .b(new_n219_), .O(new_n222_));
  OR       g0206(.a(new_n222_), .b(new_n217_), .O(new_n223_));
  OR       g0207(.a(new_n223_), .b(new_n214_), .O(new_n224_));
  OR       g0208(.a(new_n224_), .b(new_n211_), .O(new_n225_));
  AND      g0209(.a(new_n225_), .b(i_2_1_38_0), .O(new_n226_));
  OR       g0210(.a(i_2_1_70_0), .b(new_n63_), .O(new_n227_));
  AND      g0211(.a(new_n227_), .b(i_2_1_13_0), .O(new_n228_));
  AND      g0212(.a(new_n44_), .b(i_2_1_34_0), .O(new_n229_));
  NOT      g0213(.a(new_n229_), .O(new_n230_));
  OR       g0214(.a(new_n54_), .b(i_2_1_41_0), .O(new_n231_));
  OR       g0215(.a(new_n231_), .b(new_n28_), .O(new_n232_));
  NAND     g0216(.a(new_n232_), .b(new_n230_), .O(new_n233_));
  OR       g0217(.a(new_n233_), .b(new_n228_), .O(new_n234_));
  OR       g0218(.a(new_n234_), .b(new_n154_), .O(new_n235_));
  AND      g0219(.a(new_n235_), .b(new_n32_), .O(new_n236_));
  AND      g0220(.a(i_2_1_68_0), .b(i_2_1_34_0), .O(new_n237_));
  NOT      g0221(.a(new_n237_), .O(new_n238_));
  OR       g0222(.a(new_n238_), .b(new_n127_), .O(new_n239_));
  NAND     g0223(.a(new_n124_), .b(new_n220_), .O(new_n240_));
  NAND     g0224(.a(new_n240_), .b(new_n239_), .O(new_n241_));
  AND      g0225(.a(new_n241_), .b(new_n63_), .O(new_n242_));
  AND      g0226(.a(new_n39_), .b(i_2_1_34_0), .O(new_n243_));
  AND      g0227(.a(new_n73_), .b(new_n32_), .O(new_n244_));
  OR       g0228(.a(new_n244_), .b(new_n243_), .O(new_n245_));
  AND      g0229(.a(new_n245_), .b(i_2_1_49_0), .O(new_n246_));
  NOT      g0230(.a(new_n37_), .O(new_n247_));
  NAND     g0231(.a(new_n232_), .b(new_n247_), .O(new_n248_));
  AND      g0232(.a(new_n248_), .b(i_2_1_13_0), .O(new_n249_));
  OR       g0233(.a(new_n249_), .b(new_n246_), .O(new_n250_));
  OR       g0234(.a(new_n250_), .b(new_n242_), .O(new_n251_));
  OR       g0235(.a(new_n251_), .b(new_n236_), .O(new_n252_));
  OR       g0236(.a(new_n252_), .b(new_n226_), .O(new_n253_));
  AND      g0237(.a(new_n253_), .b(new_n20_), .O(new_n254_));
  NOT      g0238(.a(new_n74_), .O(new_n255_));
  OR       g0239(.a(i_2_1_135_0), .b(i_2_1_49_0), .O(new_n256_));
  OR       g0240(.a(new_n20_), .b(i_2_1_41_0), .O(new_n257_));
  OR       g0241(.a(new_n257_), .b(new_n256_), .O(new_n258_));
  NAND     g0242(.a(new_n258_), .b(new_n255_), .O(new_n259_));
  AND      g0243(.a(new_n259_), .b(new_n32_), .O(new_n260_));
  AND      g0244(.a(i_2_1_70_0), .b(i_2_1_13_0), .O(new_n261_));
  AND      g0245(.a(new_n261_), .b(new_n54_), .O(new_n262_));
  OR       g0246(.a(new_n262_), .b(new_n260_), .O(new_n263_));
  AND      g0247(.a(new_n263_), .b(i_2_1_136_0), .O(new_n264_));
  OR       g0248(.a(i_2_1_70_0), .b(i_2_1_34_0), .O(new_n265_));
  OR       g0249(.a(i_2_1_38_0), .b(i_2_1_13_0), .O(new_n266_));
  AND      g0250(.a(new_n266_), .b(new_n265_), .O(new_n267_));
  AND      g0251(.a(new_n142_), .b(i_2_1_135_0), .O(new_n268_));
  OR       g0252(.a(new_n268_), .b(new_n267_), .O(new_n269_));
  AND      g0253(.a(new_n269_), .b(new_n32_), .O(new_n270_));
  AND      g0254(.a(i_2_1_135_0), .b(new_n63_), .O(new_n271_));
  OR       g0255(.a(i_2_1_34_0), .b(i_2_1_13_0), .O(new_n272_));
  AND      g0256(.a(new_n272_), .b(i_2_1_38_0), .O(new_n273_));
  AND      g0257(.a(new_n273_), .b(new_n271_), .O(new_n274_));
  OR       g0258(.a(new_n274_), .b(new_n270_), .O(new_n275_));
  OR       g0259(.a(new_n275_), .b(new_n264_), .O(new_n276_));
  AND      g0260(.a(new_n276_), .b(i_2_1_68_0), .O(new_n277_));
  AND      g0261(.a(i_2_1_136_0), .b(i_2_1_70_0), .O(new_n278_));
  AND      g0262(.a(i_2_1_38_0), .b(i_2_1_34_0), .O(new_n279_));
  AND      g0263(.a(new_n271_), .b(new_n167_), .O(new_n280_));
  OR       g0264(.a(new_n280_), .b(new_n279_), .O(new_n281_));
  AND      g0265(.a(new_n281_), .b(new_n278_), .O(new_n282_));
  OR       g0266(.a(i_2_1_135_0), .b(i_2_1_38_0), .O(new_n283_));
  AND      g0267(.a(new_n283_), .b(new_n32_), .O(new_n284_));
  OR       g0268(.a(new_n284_), .b(new_n73_), .O(new_n285_));
  AND      g0269(.a(new_n285_), .b(new_n63_), .O(new_n286_));
  AND      g0270(.a(i_2_1_136_0), .b(i_2_1_38_0), .O(new_n287_));
  OR       g0271(.a(new_n287_), .b(new_n74_), .O(new_n288_));
  OR       g0272(.a(new_n288_), .b(new_n286_), .O(new_n289_));
  AND      g0273(.a(new_n289_), .b(new_n228_), .O(new_n290_));
  OR       g0274(.a(new_n290_), .b(new_n282_), .O(new_n291_));
  OR       g0275(.a(new_n291_), .b(new_n277_), .O(new_n292_));
  OR       g0276(.a(new_n292_), .b(new_n254_), .O(new_n293_));
  OR       g0277(.a(new_n293_), .b(new_n208_), .O(new_n294_));
  OR       g0278(.a(new_n294_), .b(new_n139_), .O(new_n295_));
  AND      g0279(.a(new_n295_), .b(i_2_1_32_0), .O(new_n296_));
  NAND     g0280(.a(new_n218_), .b(i_2_1_49_0), .O(new_n297_));
  AND      g0281(.a(new_n127_), .b(new_n93_), .O(new_n298_));
  AND      g0282(.a(new_n298_), .b(new_n297_), .O(new_n299_));
  NAND     g0283(.a(new_n128_), .b(new_n63_), .O(new_n300_));
  NAND     g0284(.a(new_n22_), .b(i_2_1_38_0), .O(new_n301_));
  NAND     g0285(.a(new_n301_), .b(new_n300_), .O(new_n302_));
  OR       g0286(.a(new_n302_), .b(new_n299_), .O(new_n303_));
  AND      g0287(.a(new_n303_), .b(new_n19_), .O(new_n304_));
  AND      g0288(.a(new_n84_), .b(new_n19_), .O(new_n305_));
  OR       g0289(.a(new_n123_), .b(i_2_1_136_0), .O(new_n306_));
  OR       g0290(.a(new_n306_), .b(new_n63_), .O(new_n307_));
  AND      g0291(.a(new_n307_), .b(new_n305_), .O(new_n308_));
  AND      g0292(.a(new_n271_), .b(i_2_1_136_0), .O(new_n309_));
  AND      g0293(.a(new_n309_), .b(new_n93_), .O(new_n310_));
  AND      g0294(.a(new_n287_), .b(new_n63_), .O(new_n311_));
  OR       g0295(.a(new_n311_), .b(new_n125_), .O(new_n312_));
  OR       g0296(.a(new_n312_), .b(new_n310_), .O(new_n313_));
  OR       g0297(.a(new_n313_), .b(new_n308_), .O(new_n314_));
  AND      g0298(.a(new_n314_), .b(i_2_1_41_0), .O(new_n315_));
  NAND     g0299(.a(new_n189_), .b(new_n53_), .O(new_n316_));
  AND      g0300(.a(new_n316_), .b(new_n82_), .O(new_n317_));
  OR       g0301(.a(new_n317_), .b(new_n315_), .O(new_n318_));
  OR       g0302(.a(new_n318_), .b(new_n304_), .O(new_n319_));
  AND      g0303(.a(new_n319_), .b(i_2_1_13_0), .O(new_n320_));
  OR       g0304(.a(new_n21_), .b(i_2_1_41_0), .O(new_n321_));
  AND      g0305(.a(new_n22_), .b(new_n63_), .O(new_n322_));
  AND      g0306(.a(new_n322_), .b(new_n321_), .O(new_n323_));
  AND      g0307(.a(i_2_1_70_0), .b(new_n63_), .O(new_n324_));
  OR       g0308(.a(new_n324_), .b(new_n32_), .O(new_n325_));
  AND      g0309(.a(new_n325_), .b(new_n127_), .O(new_n326_));
  OR       g0310(.a(i_2_1_41_0), .b(i_2_1_38_0), .O(new_n327_));
  OR       g0311(.a(i_2_1_135_0), .b(new_n32_), .O(new_n328_));
  AND      g0312(.a(new_n328_), .b(new_n327_), .O(new_n329_));
  NAND     g0313(.a(i_2_1_57_0), .b(i_2_1_54_0), .O(new_n330_));
  AND      g0314(.a(new_n330_), .b(i_2_1_13_0), .O(new_n331_));
  OR       g0315(.a(new_n331_), .b(new_n124_), .O(new_n332_));
  OR       g0316(.a(new_n332_), .b(new_n329_), .O(new_n333_));
  OR       g0317(.a(new_n333_), .b(new_n326_), .O(new_n334_));
  OR       g0318(.a(new_n334_), .b(new_n323_), .O(new_n335_));
  AND      g0319(.a(new_n335_), .b(new_n19_), .O(new_n336_));
  OR       g0320(.a(i_2_1_49_0), .b(i_2_1_46_0), .O(new_n337_));
  NOT      g0321(.a(new_n337_), .O(new_n338_));
  OR       g0322(.a(new_n338_), .b(new_n51_), .O(new_n339_));
  OR       g0323(.a(new_n339_), .b(new_n125_), .O(new_n340_));
  AND      g0324(.a(new_n340_), .b(new_n140_), .O(new_n341_));
  AND      g0325(.a(new_n63_), .b(i_2_1_41_0), .O(new_n342_));
  NOT      g0326(.a(new_n342_), .O(new_n343_));
  NAND     g0327(.a(new_n343_), .b(new_n114_), .O(new_n344_));
  AND      g0328(.a(new_n344_), .b(new_n20_), .O(new_n345_));
  AND      g0329(.a(i_2_1_49_0), .b(i_2_1_38_0), .O(new_n346_));
  AND      g0330(.a(i_2_1_135_0), .b(i_2_1_13_0), .O(new_n347_));
  OR       g0331(.a(new_n347_), .b(new_n346_), .O(new_n348_));
  AND      g0332(.a(new_n348_), .b(i_2_1_136_0), .O(new_n349_));
  OR       g0333(.a(new_n349_), .b(new_n345_), .O(new_n350_));
  OR       g0334(.a(new_n350_), .b(new_n341_), .O(new_n351_));
  NAND     g0335(.a(i_2_1_136_0), .b(i_2_1_49_0), .O(new_n352_));
  AND      g0336(.a(new_n127_), .b(i_2_1_70_0), .O(new_n353_));
  AND      g0337(.a(new_n353_), .b(new_n352_), .O(new_n354_));
  OR       g0338(.a(new_n354_), .b(new_n220_), .O(new_n355_));
  AND      g0339(.a(new_n80_), .b(i_2_1_49_0), .O(new_n356_));
  AND      g0340(.a(new_n356_), .b(new_n118_), .O(new_n357_));
  AND      g0341(.a(i_2_1_136_0), .b(i_2_1_13_0), .O(new_n358_));
  OR       g0342(.a(new_n358_), .b(i_2_1_41_0), .O(new_n359_));
  OR       g0343(.a(new_n359_), .b(new_n357_), .O(new_n360_));
  AND      g0344(.a(new_n360_), .b(new_n355_), .O(new_n361_));
  OR       g0345(.a(i_2_1_135_0), .b(i_2_1_41_0), .O(new_n362_));
  AND      g0346(.a(new_n362_), .b(new_n149_), .O(new_n363_));
  AND      g0347(.a(i_2_1_135_0), .b(i_2_1_41_0), .O(new_n364_));
  AND      g0348(.a(new_n63_), .b(i_2_1_13_0), .O(new_n365_));
  OR       g0349(.a(new_n365_), .b(new_n364_), .O(new_n366_));
  OR       g0350(.a(new_n366_), .b(new_n363_), .O(new_n367_));
  AND      g0351(.a(new_n367_), .b(new_n32_), .O(new_n368_));
  OR       g0352(.a(new_n368_), .b(new_n361_), .O(new_n369_));
  OR       g0353(.a(new_n369_), .b(new_n351_), .O(new_n370_));
  OR       g0354(.a(new_n370_), .b(new_n336_), .O(new_n371_));
  AND      g0355(.a(new_n371_), .b(i_2_1_34_0), .O(new_n372_));
  OR       g0356(.a(i_2_1_136_0), .b(i_2_1_70_0), .O(new_n373_));
  AND      g0357(.a(new_n373_), .b(i_2_1_41_0), .O(new_n374_));
  OR       g0358(.a(new_n374_), .b(new_n153_), .O(new_n375_));
  AND      g0359(.a(new_n375_), .b(new_n19_), .O(new_n376_));
  AND      g0360(.a(new_n365_), .b(i_2_1_136_0), .O(new_n377_));
  OR       g0361(.a(new_n377_), .b(new_n376_), .O(new_n378_));
  AND      g0362(.a(new_n378_), .b(i_2_1_135_0), .O(new_n379_));
  AND      g0363(.a(new_n19_), .b(i_2_1_13_0), .O(new_n380_));
  OR       g0364(.a(new_n342_), .b(new_n19_), .O(new_n381_));
  AND      g0365(.a(new_n381_), .b(new_n21_), .O(new_n382_));
  OR       g0366(.a(new_n382_), .b(new_n380_), .O(new_n383_));
  AND      g0367(.a(new_n383_), .b(new_n93_), .O(new_n384_));
  OR       g0368(.a(new_n380_), .b(new_n199_), .O(new_n385_));
  AND      g0369(.a(new_n385_), .b(i_2_1_38_0), .O(new_n386_));
  AND      g0370(.a(i_2_1_41_0), .b(i_2_1_13_0), .O(new_n387_));
  AND      g0371(.a(new_n387_), .b(new_n84_), .O(new_n388_));
  OR       g0372(.a(i_2_1_136_0), .b(new_n20_), .O(new_n389_));
  AND      g0373(.a(new_n389_), .b(new_n63_), .O(new_n390_));
  AND      g0374(.a(new_n390_), .b(new_n305_), .O(new_n391_));
  OR       g0375(.a(new_n391_), .b(new_n388_), .O(new_n392_));
  OR       g0376(.a(new_n392_), .b(new_n386_), .O(new_n393_));
  OR       g0377(.a(new_n393_), .b(new_n384_), .O(new_n394_));
  OR       g0378(.a(new_n394_), .b(new_n379_), .O(new_n395_));
  AND      g0379(.a(new_n395_), .b(new_n32_), .O(new_n396_));
  AND      g0380(.a(i_2_1_70_0), .b(new_n19_), .O(new_n397_));
  AND      g0381(.a(new_n397_), .b(new_n199_), .O(new_n398_));
  OR       g0382(.a(new_n54_), .b(i_2_1_57_0), .O(new_n399_));
  OR       g0383(.a(new_n399_), .b(new_n27_), .O(new_n400_));
  NAND     g0384(.a(new_n397_), .b(new_n65_), .O(new_n401_));
  NAND     g0385(.a(new_n401_), .b(new_n400_), .O(new_n402_));
  OR       g0386(.a(i_2_1_70_0), .b(new_n19_), .O(new_n403_));
  AND      g0387(.a(new_n403_), .b(new_n389_), .O(new_n404_));
  AND      g0388(.a(new_n404_), .b(i_2_1_41_0), .O(new_n405_));
  AND      g0389(.a(new_n405_), .b(new_n402_), .O(new_n406_));
  OR       g0390(.a(new_n406_), .b(new_n398_), .O(new_n407_));
  AND      g0391(.a(new_n407_), .b(new_n63_), .O(new_n408_));
  OR       g0392(.a(new_n389_), .b(new_n63_), .O(new_n409_));
  AND      g0393(.a(new_n409_), .b(i_2_1_70_0), .O(new_n410_));
  OR       g0394(.a(new_n410_), .b(i_2_1_41_0), .O(new_n411_));
  AND      g0395(.a(i_2_1_136_0), .b(new_n53_), .O(new_n412_));
  OR       g0396(.a(i_2_1_135_0), .b(i_2_1_46_0), .O(new_n413_));
  NOT      g0397(.a(new_n413_), .O(new_n414_));
  OR       g0398(.a(new_n414_), .b(new_n412_), .O(new_n415_));
  NAND     g0399(.a(new_n415_), .b(i_2_1_49_0), .O(new_n416_));
  AND      g0400(.a(new_n93_), .b(i_2_1_136_0), .O(new_n417_));
  OR       g0401(.a(new_n417_), .b(new_n19_), .O(new_n418_));
  AND      g0402(.a(new_n418_), .b(new_n416_), .O(new_n419_));
  OR       g0403(.a(new_n33_), .b(i_2_1_136_0), .O(new_n420_));
  AND      g0404(.a(new_n420_), .b(i_2_1_38_0), .O(new_n421_));
  OR       g0405(.a(new_n404_), .b(i_2_1_135_0), .O(new_n422_));
  AND      g0406(.a(new_n422_), .b(new_n421_), .O(new_n423_));
  AND      g0407(.a(new_n423_), .b(new_n419_), .O(new_n424_));
  AND      g0408(.a(new_n424_), .b(new_n411_), .O(new_n425_));
  OR       g0409(.a(new_n425_), .b(new_n408_), .O(new_n426_));
  OR       g0410(.a(new_n426_), .b(new_n396_), .O(new_n427_));
  OR       g0411(.a(new_n427_), .b(new_n372_), .O(new_n428_));
  OR       g0412(.a(new_n428_), .b(new_n320_), .O(new_n429_));
  AND      g0413(.a(new_n429_), .b(i_2_1_68_0), .O(new_n430_));
  AND      g0414(.a(i_2_1_136_0), .b(i_2_1_41_0), .O(new_n431_));
  OR       g0415(.a(new_n431_), .b(new_n397_), .O(new_n432_));
  AND      g0416(.a(new_n432_), .b(new_n20_), .O(new_n433_));
  OR       g0417(.a(new_n433_), .b(new_n123_), .O(new_n434_));
  AND      g0418(.a(new_n434_), .b(new_n32_), .O(new_n435_));
  OR       g0419(.a(i_2_1_57_0), .b(i_2_1_46_0), .O(new_n436_));
  NAND     g0420(.a(new_n436_), .b(i_2_1_136_0), .O(new_n437_));
  AND      g0421(.a(i_2_1_70_0), .b(i_2_1_41_0), .O(new_n438_));
  OR       g0422(.a(new_n438_), .b(i_2_1_136_0), .O(new_n439_));
  AND      g0423(.a(new_n193_), .b(i_2_1_54_0), .O(new_n440_));
  AND      g0424(.a(new_n440_), .b(new_n439_), .O(new_n441_));
  AND      g0425(.a(new_n441_), .b(new_n437_), .O(new_n442_));
  OR       g0426(.a(new_n124_), .b(new_n80_), .O(new_n443_));
  AND      g0427(.a(new_n443_), .b(i_2_1_13_0), .O(new_n444_));
  AND      g0428(.a(new_n19_), .b(i_2_1_41_0), .O(new_n445_));
  OR       g0429(.a(new_n54_), .b(i_2_1_70_0), .O(new_n446_));
  AND      g0430(.a(new_n446_), .b(new_n445_), .O(new_n447_));
  NOT      g0431(.a(new_n111_), .O(new_n448_));
  OR       g0432(.a(new_n397_), .b(new_n448_), .O(new_n449_));
  AND      g0433(.a(new_n449_), .b(i_2_1_34_0), .O(new_n450_));
  OR       g0434(.a(new_n450_), .b(new_n447_), .O(new_n451_));
  OR       g0435(.a(new_n451_), .b(new_n444_), .O(new_n452_));
  OR       g0436(.a(new_n452_), .b(new_n442_), .O(new_n453_));
  OR       g0437(.a(new_n453_), .b(new_n435_), .O(new_n454_));
  AND      g0438(.a(new_n454_), .b(new_n63_), .O(new_n455_));
  AND      g0439(.a(new_n438_), .b(i_2_1_136_0), .O(new_n456_));
  OR       g0440(.a(new_n456_), .b(new_n64_), .O(new_n457_));
  AND      g0441(.a(new_n457_), .b(i_2_1_13_0), .O(new_n458_));
  NOT      g0442(.a(new_n431_), .O(new_n459_));
  NAND     g0443(.a(new_n459_), .b(new_n111_), .O(new_n460_));
  AND      g0444(.a(new_n460_), .b(new_n20_), .O(new_n461_));
  AND      g0445(.a(new_n178_), .b(new_n33_), .O(new_n462_));
  AND      g0446(.a(i_2_1_70_0), .b(new_n32_), .O(new_n463_));
  AND      g0447(.a(new_n463_), .b(i_2_1_34_0), .O(new_n464_));
  OR       g0448(.a(new_n464_), .b(i_2_1_46_0), .O(new_n465_));
  OR       g0449(.a(new_n465_), .b(new_n462_), .O(new_n466_));
  OR       g0450(.a(new_n466_), .b(new_n461_), .O(new_n467_));
  OR       g0451(.a(new_n467_), .b(new_n458_), .O(new_n468_));
  NAND     g0452(.a(i_2_1_54_0), .b(i_2_1_49_0), .O(new_n469_));
  AND      g0453(.a(i_2_1_34_0), .b(i_2_1_13_0), .O(new_n470_));
  NOT      g0454(.a(new_n470_), .O(new_n471_));
  OR       g0455(.a(new_n471_), .b(new_n469_), .O(new_n472_));
  AND      g0456(.a(new_n112_), .b(i_2_1_46_0), .O(new_n473_));
  NAND     g0457(.a(new_n473_), .b(new_n472_), .O(new_n474_));
  AND      g0458(.a(new_n474_), .b(new_n468_), .O(new_n475_));
  NAND     g0459(.a(new_n306_), .b(new_n32_), .O(new_n476_));
  OR       g0460(.a(new_n164_), .b(i_2_1_57_0), .O(new_n477_));
  NAND     g0461(.a(new_n477_), .b(new_n476_), .O(new_n478_));
  AND      g0462(.a(new_n478_), .b(i_2_1_13_0), .O(new_n479_));
  AND      g0463(.a(new_n403_), .b(i_2_1_41_0), .O(new_n480_));
  NAND     g0464(.a(new_n362_), .b(i_2_1_13_0), .O(new_n481_));
  NAND     g0465(.a(new_n481_), .b(new_n400_), .O(new_n482_));
  OR       g0466(.a(new_n482_), .b(new_n480_), .O(new_n483_));
  AND      g0467(.a(new_n483_), .b(i_2_1_34_0), .O(new_n484_));
  OR       g0468(.a(new_n484_), .b(new_n479_), .O(new_n485_));
  OR       g0469(.a(new_n485_), .b(new_n475_), .O(new_n486_));
  OR       g0470(.a(new_n486_), .b(new_n455_), .O(new_n487_));
  AND      g0471(.a(new_n487_), .b(i_2_1_38_0), .O(new_n488_));
  AND      g0472(.a(i_2_1_135_0), .b(new_n19_), .O(new_n489_));
  AND      g0473(.a(new_n489_), .b(i_2_1_34_0), .O(new_n490_));
  OR       g0474(.a(new_n490_), .b(new_n148_), .O(new_n491_));
  AND      g0475(.a(new_n491_), .b(i_2_1_70_0), .O(new_n492_));
  OR       g0476(.a(i_2_1_135_0), .b(new_n19_), .O(new_n493_));
  NAND     g0477(.a(new_n493_), .b(i_2_1_34_0), .O(new_n494_));
  OR       g0478(.a(i_2_1_46_0), .b(i_2_1_38_0), .O(new_n495_));
  OR       g0479(.a(new_n495_), .b(new_n27_), .O(new_n496_));
  NAND     g0480(.a(new_n496_), .b(new_n494_), .O(new_n497_));
  AND      g0481(.a(new_n497_), .b(new_n63_), .O(new_n498_));
  OR       g0482(.a(new_n431_), .b(new_n271_), .O(new_n499_));
  AND      g0483(.a(new_n499_), .b(i_2_1_13_0), .O(new_n500_));
  OR       g0484(.a(new_n500_), .b(new_n480_), .O(new_n501_));
  OR       g0485(.a(new_n501_), .b(new_n498_), .O(new_n502_));
  OR       g0486(.a(new_n502_), .b(new_n492_), .O(new_n503_));
  AND      g0487(.a(new_n503_), .b(new_n32_), .O(new_n504_));
  AND      g0488(.a(new_n387_), .b(new_n32_), .O(new_n505_));
  AND      g0489(.a(new_n212_), .b(i_2_1_70_0), .O(new_n506_));
  OR       g0490(.a(new_n506_), .b(new_n505_), .O(new_n507_));
  AND      g0491(.a(new_n507_), .b(new_n54_), .O(new_n508_));
  AND      g0492(.a(new_n347_), .b(i_2_1_34_0), .O(new_n509_));
  AND      g0493(.a(new_n321_), .b(new_n261_), .O(new_n510_));
  OR       g0494(.a(new_n510_), .b(new_n509_), .O(new_n511_));
  OR       g0495(.a(new_n511_), .b(new_n508_), .O(new_n512_));
  OR       g0496(.a(new_n512_), .b(new_n504_), .O(new_n513_));
  AND      g0497(.a(new_n513_), .b(new_n20_), .O(new_n514_));
  OR       g0498(.a(new_n489_), .b(i_2_1_136_0), .O(new_n515_));
  OR       g0499(.a(new_n463_), .b(i_2_1_13_0), .O(new_n516_));
  AND      g0500(.a(new_n516_), .b(new_n515_), .O(new_n517_));
  OR       g0501(.a(new_n278_), .b(new_n32_), .O(new_n518_));
  AND      g0502(.a(new_n518_), .b(new_n445_), .O(new_n519_));
  OR       g0503(.a(new_n519_), .b(new_n517_), .O(new_n520_));
  AND      g0504(.a(new_n520_), .b(new_n63_), .O(new_n521_));
  OR       g0505(.a(new_n397_), .b(new_n21_), .O(new_n522_));
  AND      g0506(.a(new_n522_), .b(i_2_1_13_0), .O(new_n523_));
  AND      g0507(.a(i_2_1_49_0), .b(i_2_1_41_0), .O(new_n524_));
  OR       g0508(.a(new_n524_), .b(i_2_1_136_0), .O(new_n525_));
  AND      g0509(.a(new_n525_), .b(new_n123_), .O(new_n526_));
  OR       g0510(.a(new_n526_), .b(new_n523_), .O(new_n527_));
  AND      g0511(.a(new_n527_), .b(new_n32_), .O(new_n528_));
  OR       g0512(.a(new_n528_), .b(new_n521_), .O(new_n529_));
  AND      g0513(.a(new_n529_), .b(i_2_1_34_0), .O(new_n530_));
  NOT      g0514(.a(i_2_1_13_0), .O(new_n531_));
  AND      g0515(.a(i_2_1_41_0), .b(i_2_1_38_0), .O(new_n532_));
  NOT      g0516(.a(new_n532_), .O(new_n533_));
  OR       g0517(.a(new_n533_), .b(new_n86_), .O(new_n534_));
  AND      g0518(.a(i_2_1_34_0), .b(i_2_1_32_0), .O(new_n535_));
  NOT      g0519(.a(new_n535_), .O(new_n536_));
  OR       g0520(.a(new_n256_), .b(new_n193_), .O(new_n537_));
  OR       g0521(.a(new_n537_), .b(new_n536_), .O(new_n538_));
  NAND     g0522(.a(new_n538_), .b(new_n534_), .O(new_n539_));
  AND      g0523(.a(new_n539_), .b(new_n531_), .O(new_n540_));
  OR       g0524(.a(new_n278_), .b(new_n82_), .O(new_n541_));
  AND      g0525(.a(new_n541_), .b(new_n19_), .O(new_n542_));
  OR       g0526(.a(new_n542_), .b(new_n278_), .O(new_n543_));
  NAND     g0527(.a(new_n535_), .b(new_n32_), .O(new_n544_));
  OR       g0528(.a(i_2_1_32_0), .b(new_n531_), .O(new_n545_));
  OR       g0529(.a(new_n545_), .b(i_2_1_57_0), .O(new_n546_));
  NAND     g0530(.a(new_n546_), .b(new_n544_), .O(new_n547_));
  NAND     g0531(.a(new_n547_), .b(new_n543_), .O(new_n548_));
  AND      g0532(.a(i_2_1_136_0), .b(new_n19_), .O(new_n549_));
  NAND     g0533(.a(new_n549_), .b(i_2_1_41_0), .O(new_n550_));
  AND      g0534(.a(new_n550_), .b(i_2_1_54_0), .O(new_n551_));
  OR       g0535(.a(new_n271_), .b(new_n178_), .O(new_n552_));
  NAND     g0536(.a(new_n552_), .b(new_n261_), .O(new_n553_));
  OR       g0537(.a(new_n553_), .b(new_n551_), .O(new_n554_));
  NAND     g0538(.a(new_n554_), .b(new_n548_), .O(new_n555_));
  OR       g0539(.a(new_n555_), .b(new_n540_), .O(new_n556_));
  OR       g0540(.a(new_n556_), .b(new_n530_), .O(new_n557_));
  OR       g0541(.a(new_n557_), .b(new_n514_), .O(new_n558_));
  OR       g0542(.a(new_n558_), .b(new_n488_), .O(new_n559_));
  OR       g0543(.a(new_n559_), .b(new_n430_), .O(new_n560_));
  OR       g0544(.a(new_n560_), .b(new_n296_), .O(new_n561_));
  AND      g0545(.a(new_n561_), .b(new_n18_), .O(new_n562_));
  OR       g0546(.a(new_n337_), .b(new_n18_), .O(new_n563_));
  OR       g0547(.a(new_n563_), .b(i_2_1_70_0), .O(new_n564_));
  NAND     g0548(.a(new_n564_), .b(new_n218_), .O(new_n565_));
  AND      g0549(.a(new_n565_), .b(new_n220_), .O(new_n566_));
  AND      g0550(.a(i_2_1_68_0), .b(i_2_1_41_0), .O(new_n567_));
  OR       g0551(.a(new_n567_), .b(i_2_1_70_0), .O(new_n568_));
  AND      g0552(.a(new_n568_), .b(i_2_1_135_0), .O(new_n569_));
  OR       g0553(.a(new_n237_), .b(i_2_1_136_0), .O(new_n570_));
  AND      g0554(.a(new_n570_), .b(new_n63_), .O(new_n571_));
  OR       g0555(.a(new_n571_), .b(new_n569_), .O(new_n572_));
  AND      g0556(.a(i_2_1_70_0), .b(i_2_1_51_0), .O(new_n573_));
  OR       g0557(.a(new_n25_), .b(i_2_1_46_0), .O(new_n574_));
  NOT      g0558(.a(new_n574_), .O(new_n575_));
  OR       g0559(.a(new_n575_), .b(new_n573_), .O(new_n576_));
  AND      g0560(.a(new_n576_), .b(i_2_1_34_0), .O(new_n577_));
  OR       g0561(.a(new_n279_), .b(new_n51_), .O(new_n578_));
  AND      g0562(.a(new_n578_), .b(i_2_1_68_0), .O(new_n579_));
  OR       g0563(.a(new_n532_), .b(i_2_1_70_0), .O(new_n580_));
  AND      g0564(.a(new_n580_), .b(new_n327_), .O(new_n581_));
  OR       g0565(.a(new_n581_), .b(new_n579_), .O(new_n582_));
  OR       g0566(.a(new_n582_), .b(new_n577_), .O(new_n583_));
  OR       g0567(.a(new_n583_), .b(new_n572_), .O(new_n584_));
  OR       g0568(.a(new_n584_), .b(new_n566_), .O(new_n585_));
  AND      g0569(.a(new_n585_), .b(i_2_1_13_0), .O(new_n586_));
  AND      g0570(.a(new_n149_), .b(i_2_1_34_0), .O(new_n587_));
  AND      g0571(.a(i_2_1_51_0), .b(new_n19_), .O(new_n588_));
  AND      g0572(.a(new_n588_), .b(new_n169_), .O(new_n589_));
  OR       g0573(.a(new_n589_), .b(new_n549_), .O(new_n590_));
  OR       g0574(.a(new_n590_), .b(new_n421_), .O(new_n591_));
  OR       g0575(.a(new_n591_), .b(new_n587_), .O(new_n592_));
  AND      g0576(.a(new_n592_), .b(i_2_1_41_0), .O(new_n593_));
  NAND     g0577(.a(i_2_1_49_0), .b(i_2_1_46_0), .O(new_n594_));
  AND      g0578(.a(new_n594_), .b(i_2_1_34_0), .O(new_n595_));
  OR       g0579(.a(new_n338_), .b(new_n68_), .O(new_n596_));
  AND      g0580(.a(new_n596_), .b(new_n595_), .O(new_n597_));
  AND      g0581(.a(new_n338_), .b(i_2_1_38_0), .O(new_n598_));
  OR       g0582(.a(new_n324_), .b(new_n279_), .O(new_n599_));
  AND      g0583(.a(new_n599_), .b(i_2_1_136_0), .O(new_n600_));
  OR       g0584(.a(new_n600_), .b(new_n598_), .O(new_n601_));
  OR       g0585(.a(new_n601_), .b(new_n597_), .O(new_n602_));
  OR       g0586(.a(new_n602_), .b(new_n593_), .O(new_n603_));
  AND      g0587(.a(new_n603_), .b(i_2_1_68_0), .O(new_n604_));
  AND      g0588(.a(new_n342_), .b(new_n278_), .O(new_n605_));
  AND      g0589(.a(new_n141_), .b(i_2_1_136_0), .O(new_n606_));
  OR       g0590(.a(new_n148_), .b(i_2_1_34_0), .O(new_n607_));
  AND      g0591(.a(new_n607_), .b(i_2_1_38_0), .O(new_n608_));
  AND      g0592(.a(new_n141_), .b(i_2_1_41_0), .O(new_n609_));
  OR       g0593(.a(new_n609_), .b(new_n608_), .O(new_n610_));
  AND      g0594(.a(new_n610_), .b(i_2_1_70_0), .O(new_n611_));
  OR       g0595(.a(new_n611_), .b(new_n606_), .O(new_n612_));
  AND      g0596(.a(new_n612_), .b(new_n19_), .O(new_n613_));
  OR       g0597(.a(new_n613_), .b(new_n605_), .O(new_n614_));
  OR       g0598(.a(new_n614_), .b(new_n604_), .O(new_n615_));
  OR       g0599(.a(new_n615_), .b(new_n586_), .O(new_n616_));
  OR       g0600(.a(new_n18_), .b(i_2_1_41_0), .O(new_n617_));
  NOT      g0601(.a(new_n617_), .O(new_n618_));
  OR       g0602(.a(new_n94_), .b(new_n53_), .O(new_n619_));
  NAND     g0603(.a(new_n619_), .b(new_n255_), .O(new_n620_));
  AND      g0604(.a(new_n620_), .b(new_n618_), .O(new_n621_));
  OR       g0605(.a(new_n621_), .b(new_n237_), .O(new_n622_));
  AND      g0606(.a(new_n622_), .b(i_2_1_136_0), .O(new_n623_));
  NOT      g0607(.a(new_n438_), .O(new_n624_));
  NAND     g0608(.a(new_n380_), .b(i_2_1_51_0), .O(new_n625_));
  OR       g0609(.a(new_n625_), .b(i_2_1_135_0), .O(new_n626_));
  NAND     g0610(.a(new_n626_), .b(new_n624_), .O(new_n627_));
  AND      g0611(.a(new_n627_), .b(new_n102_), .O(new_n628_));
  AND      g0612(.a(new_n227_), .b(new_n74_), .O(new_n629_));
  OR       g0613(.a(new_n365_), .b(new_n237_), .O(new_n630_));
  AND      g0614(.a(new_n630_), .b(i_2_1_41_0), .O(new_n631_));
  OR       g0615(.a(new_n631_), .b(new_n629_), .O(new_n632_));
  OR       g0616(.a(new_n632_), .b(new_n628_), .O(new_n633_));
  OR       g0617(.a(new_n633_), .b(new_n623_), .O(new_n634_));
  AND      g0618(.a(i_2_1_46_0), .b(i_2_1_13_0), .O(new_n635_));
  OR       g0619(.a(i_2_1_68_0), .b(new_n19_), .O(new_n636_));
  AND      g0620(.a(new_n493_), .b(i_2_1_68_0), .O(new_n637_));
  OR       g0621(.a(i_2_1_41_0), .b(i_2_1_34_0), .O(new_n638_));
  OR       g0622(.a(new_n638_), .b(new_n324_), .O(new_n639_));
  OR       g0623(.a(new_n639_), .b(new_n637_), .O(new_n640_));
  AND      g0624(.a(new_n640_), .b(new_n636_), .O(new_n641_));
  OR       g0625(.a(new_n641_), .b(new_n635_), .O(new_n642_));
  AND      g0626(.a(new_n642_), .b(i_2_1_38_0), .O(new_n643_));
  OR       g0627(.a(new_n19_), .b(i_2_1_13_0), .O(new_n644_));
  AND      g0628(.a(new_n644_), .b(i_2_1_34_0), .O(new_n645_));
  OR       g0629(.a(new_n645_), .b(new_n347_), .O(new_n646_));
  OR       g0630(.a(new_n646_), .b(new_n311_), .O(new_n647_));
  OR       g0631(.a(new_n647_), .b(new_n382_), .O(new_n648_));
  AND      g0632(.a(new_n648_), .b(i_2_1_68_0), .O(new_n649_));
  OR       g0633(.a(new_n649_), .b(new_n643_), .O(new_n650_));
  OR       g0634(.a(new_n650_), .b(new_n634_), .O(new_n651_));
  AND      g0635(.a(new_n651_), .b(new_n20_), .O(new_n652_));
  OR       g0636(.a(new_n374_), .b(new_n63_), .O(new_n653_));
  OR       g0637(.a(new_n39_), .b(i_2_1_41_0), .O(new_n654_));
  OR       g0638(.a(new_n654_), .b(new_n573_), .O(new_n655_));
  OR       g0639(.a(new_n44_), .b(new_n19_), .O(new_n656_));
  AND      g0640(.a(new_n656_), .b(new_n655_), .O(new_n657_));
  AND      g0641(.a(new_n657_), .b(new_n653_), .O(new_n658_));
  OR       g0642(.a(new_n532_), .b(new_n278_), .O(new_n659_));
  AND      g0643(.a(i_2_1_68_0), .b(i_2_1_38_0), .O(new_n660_));
  NOT      g0644(.a(new_n660_), .O(new_n661_));
  NAND     g0645(.a(new_n661_), .b(new_n574_), .O(new_n662_));
  OR       g0646(.a(new_n662_), .b(new_n659_), .O(new_n663_));
  OR       g0647(.a(new_n663_), .b(new_n658_), .O(new_n664_));
  AND      g0648(.a(new_n664_), .b(i_2_1_34_0), .O(new_n665_));
  AND      g0649(.a(new_n68_), .b(i_2_1_136_0), .O(new_n666_));
  OR       g0650(.a(new_n666_), .b(new_n324_), .O(new_n667_));
  AND      g0651(.a(new_n667_), .b(i_2_1_68_0), .O(new_n668_));
  AND      g0652(.a(new_n148_), .b(i_2_1_68_0), .O(new_n669_));
  OR       g0653(.a(new_n73_), .b(i_2_1_46_0), .O(new_n670_));
  OR       g0654(.a(new_n670_), .b(new_n669_), .O(new_n671_));
  OR       g0655(.a(i_2_1_70_0), .b(new_n102_), .O(new_n672_));
  OR       g0656(.a(new_n672_), .b(new_n343_), .O(new_n673_));
  NOT      g0657(.a(new_n278_), .O(new_n674_));
  AND      g0658(.a(new_n674_), .b(i_2_1_46_0), .O(new_n675_));
  NAND     g0659(.a(new_n675_), .b(new_n673_), .O(new_n676_));
  AND      g0660(.a(new_n676_), .b(new_n671_), .O(new_n677_));
  OR       g0661(.a(new_n677_), .b(new_n668_), .O(new_n678_));
  OR       g0662(.a(new_n678_), .b(new_n665_), .O(new_n679_));
  AND      g0663(.a(new_n679_), .b(i_2_1_135_0), .O(new_n680_));
  OR       g0664(.a(new_n680_), .b(new_n652_), .O(new_n681_));
  OR       g0665(.a(new_n681_), .b(new_n616_), .O(new_n682_));
  AND      g0666(.a(new_n682_), .b(i_2_1_32_0), .O(new_n683_));
  OR       g0667(.a(new_n271_), .b(i_2_1_41_0), .O(new_n684_));
  AND      g0668(.a(new_n684_), .b(i_2_1_38_0), .O(new_n685_));
  AND      g0669(.a(new_n165_), .b(i_2_1_13_0), .O(new_n686_));
  OR       g0670(.a(new_n686_), .b(new_n347_), .O(new_n687_));
  OR       g0671(.a(new_n687_), .b(new_n685_), .O(new_n688_));
  OR       g0672(.a(new_n688_), .b(new_n323_), .O(new_n689_));
  AND      g0673(.a(new_n689_), .b(new_n19_), .O(new_n690_));
  AND      g0674(.a(new_n84_), .b(i_2_1_41_0), .O(new_n691_));
  OR       g0675(.a(new_n347_), .b(new_n309_), .O(new_n692_));
  OR       g0676(.a(new_n692_), .b(new_n691_), .O(new_n693_));
  NAND     g0677(.a(new_n337_), .b(new_n102_), .O(new_n694_));
  OR       g0678(.a(new_n96_), .b(new_n19_), .O(new_n695_));
  AND      g0679(.a(new_n695_), .b(new_n694_), .O(new_n696_));
  OR       g0680(.a(i_2_1_70_0), .b(i_2_1_13_0), .O(new_n697_));
  OR       g0681(.a(new_n63_), .b(i_2_1_38_0), .O(new_n698_));
  OR       g0682(.a(new_n698_), .b(new_n19_), .O(new_n699_));
  AND      g0683(.a(new_n699_), .b(new_n697_), .O(new_n700_));
  OR       g0684(.a(new_n700_), .b(new_n696_), .O(new_n701_));
  OR       g0685(.a(new_n701_), .b(new_n693_), .O(new_n702_));
  AND      g0686(.a(new_n702_), .b(i_2_1_34_0), .O(new_n703_));
  NAND     g0687(.a(new_n347_), .b(i_2_1_136_0), .O(new_n704_));
  OR       g0688(.a(new_n532_), .b(new_n175_), .O(new_n705_));
  NAND     g0689(.a(new_n705_), .b(i_2_1_70_0), .O(new_n706_));
  NAND     g0690(.a(new_n706_), .b(new_n704_), .O(new_n707_));
  AND      g0691(.a(new_n707_), .b(new_n63_), .O(new_n708_));
  AND      g0692(.a(i_2_1_38_0), .b(i_2_1_13_0), .O(new_n709_));
  OR       g0693(.a(new_n709_), .b(new_n21_), .O(new_n710_));
  AND      g0694(.a(new_n710_), .b(new_n82_), .O(new_n711_));
  AND      g0695(.a(new_n127_), .b(i_2_1_41_0), .O(new_n712_));
  OR       g0696(.a(new_n266_), .b(new_n123_), .O(new_n713_));
  AND      g0697(.a(new_n713_), .b(new_n712_), .O(new_n714_));
  OR       g0698(.a(new_n714_), .b(new_n711_), .O(new_n715_));
  OR       g0699(.a(new_n715_), .b(new_n708_), .O(new_n716_));
  OR       g0700(.a(new_n716_), .b(new_n703_), .O(new_n717_));
  OR       g0701(.a(new_n717_), .b(new_n690_), .O(new_n718_));
  AND      g0702(.a(new_n718_), .b(i_2_1_68_0), .O(new_n719_));
  OR       g0703(.a(new_n397_), .b(i_2_1_34_0), .O(new_n720_));
  AND      g0704(.a(new_n720_), .b(i_2_1_41_0), .O(new_n721_));
  OR       g0705(.a(new_n549_), .b(i_2_1_135_0), .O(new_n722_));
  AND      g0706(.a(new_n722_), .b(i_2_1_70_0), .O(new_n723_));
  OR       g0707(.a(new_n723_), .b(new_n721_), .O(new_n724_));
  AND      g0708(.a(new_n724_), .b(new_n63_), .O(new_n725_));
  NAND     g0709(.a(new_n697_), .b(i_2_1_34_0), .O(new_n726_));
  OR       g0710(.a(new_n27_), .b(i_2_1_41_0), .O(new_n727_));
  OR       g0711(.a(new_n727_), .b(new_n54_), .O(new_n728_));
  NAND     g0712(.a(new_n728_), .b(new_n726_), .O(new_n729_));
  AND      g0713(.a(new_n729_), .b(new_n19_), .O(new_n730_));
  OR       g0714(.a(new_n730_), .b(new_n686_), .O(new_n731_));
  OR       g0715(.a(new_n731_), .b(new_n725_), .O(new_n732_));
  AND      g0716(.a(new_n732_), .b(i_2_1_38_0), .O(new_n733_));
  AND      g0717(.a(new_n638_), .b(i_2_1_13_0), .O(new_n734_));
  OR       g0718(.a(new_n342_), .b(new_n74_), .O(new_n735_));
  AND      g0719(.a(new_n735_), .b(i_2_1_136_0), .O(new_n736_));
  OR       g0720(.a(new_n736_), .b(new_n734_), .O(new_n737_));
  AND      g0721(.a(new_n737_), .b(i_2_1_70_0), .O(new_n738_));
  NOT      g0722(.a(new_n265_), .O(new_n739_));
  AND      g0723(.a(new_n365_), .b(new_n739_), .O(new_n740_));
  AND      g0724(.a(i_2_1_41_0), .b(i_2_1_34_0), .O(new_n741_));
  AND      g0725(.a(new_n741_), .b(i_2_1_136_0), .O(new_n742_));
  OR       g0726(.a(new_n742_), .b(new_n740_), .O(new_n743_));
  AND      g0727(.a(new_n743_), .b(new_n19_), .O(new_n744_));
  OR       g0728(.a(new_n741_), .b(new_n397_), .O(new_n745_));
  NAND     g0729(.a(new_n661_), .b(new_n29_), .O(new_n746_));
  AND      g0730(.a(new_n746_), .b(new_n745_), .O(new_n747_));
  AND      g0731(.a(new_n470_), .b(i_2_1_136_0), .O(new_n748_));
  OR       g0732(.a(new_n709_), .b(new_n74_), .O(new_n749_));
  AND      g0733(.a(new_n27_), .b(i_2_1_41_0), .O(new_n750_));
  OR       g0734(.a(new_n750_), .b(new_n575_), .O(new_n751_));
  AND      g0735(.a(new_n751_), .b(new_n749_), .O(new_n752_));
  OR       g0736(.a(new_n752_), .b(new_n748_), .O(new_n753_));
  OR       g0737(.a(new_n753_), .b(new_n747_), .O(new_n754_));
  OR       g0738(.a(new_n754_), .b(new_n744_), .O(new_n755_));
  OR       g0739(.a(new_n755_), .b(new_n738_), .O(new_n756_));
  OR       g0740(.a(new_n756_), .b(new_n733_), .O(new_n757_));
  OR       g0741(.a(new_n757_), .b(new_n719_), .O(new_n758_));
  AND      g0742(.a(new_n758_), .b(new_n20_), .O(new_n759_));
  AND      g0743(.a(new_n431_), .b(i_2_1_135_0), .O(new_n760_));
  OR       g0744(.a(new_n760_), .b(new_n103_), .O(new_n761_));
  OR       g0745(.a(new_n63_), .b(i_2_1_41_0), .O(new_n762_));
  AND      g0746(.a(new_n762_), .b(new_n44_), .O(new_n763_));
  AND      g0747(.a(new_n373_), .b(i_2_1_68_0), .O(new_n764_));
  OR       g0748(.a(new_n764_), .b(new_n763_), .O(new_n765_));
  OR       g0749(.a(new_n765_), .b(new_n761_), .O(new_n766_));
  AND      g0750(.a(new_n766_), .b(i_2_1_34_0), .O(new_n767_));
  OR       g0751(.a(new_n26_), .b(new_n53_), .O(new_n768_));
  NAND     g0752(.a(new_n768_), .b(new_n459_), .O(new_n769_));
  AND      g0753(.a(new_n769_), .b(new_n44_), .O(new_n770_));
  OR       g0754(.a(new_n770_), .b(new_n767_), .O(new_n771_));
  AND      g0755(.a(new_n771_), .b(new_n19_), .O(new_n772_));
  AND      g0756(.a(new_n192_), .b(new_n21_), .O(new_n773_));
  AND      g0757(.a(new_n438_), .b(new_n209_), .O(new_n774_));
  OR       g0758(.a(new_n774_), .b(new_n773_), .O(new_n775_));
  AND      g0759(.a(new_n775_), .b(new_n155_), .O(new_n776_));
  OR       g0760(.a(new_n364_), .b(i_2_1_136_0), .O(new_n777_));
  AND      g0761(.a(new_n777_), .b(new_n37_), .O(new_n778_));
  NAND     g0762(.a(new_n549_), .b(new_n123_), .O(new_n779_));
  NOT      g0763(.a(new_n387_), .O(new_n780_));
  OR       g0764(.a(i_2_1_136_0), .b(new_n18_), .O(new_n781_));
  OR       g0765(.a(new_n781_), .b(new_n780_), .O(new_n782_));
  NAND     g0766(.a(new_n782_), .b(new_n779_), .O(new_n783_));
  AND      g0767(.a(new_n783_), .b(i_2_1_49_0), .O(new_n784_));
  OR       g0768(.a(new_n784_), .b(new_n778_), .O(new_n785_));
  OR       g0769(.a(new_n785_), .b(new_n776_), .O(new_n786_));
  OR       g0770(.a(new_n786_), .b(new_n772_), .O(new_n787_));
  AND      g0771(.a(new_n297_), .b(i_2_1_41_0), .O(new_n788_));
  OR       g0772(.a(new_n788_), .b(new_n123_), .O(new_n789_));
  AND      g0773(.a(new_n789_), .b(i_2_1_68_0), .O(new_n790_));
  AND      g0774(.a(new_n324_), .b(new_n54_), .O(new_n791_));
  OR       g0775(.a(new_n791_), .b(new_n790_), .O(new_n792_));
  AND      g0776(.a(new_n792_), .b(i_2_1_34_0), .O(new_n793_));
  OR       g0777(.a(new_n21_), .b(i_2_1_34_0), .O(new_n794_));
  OR       g0778(.a(new_n794_), .b(new_n489_), .O(new_n795_));
  AND      g0779(.a(new_n795_), .b(new_n637_), .O(new_n796_));
  AND      g0780(.a(new_n19_), .b(i_2_1_34_0), .O(new_n797_));
  OR       g0781(.a(new_n797_), .b(i_2_1_68_0), .O(new_n798_));
  AND      g0782(.a(new_n798_), .b(i_2_1_70_0), .O(new_n799_));
  AND      g0783(.a(new_n175_), .b(i_2_1_41_0), .O(new_n800_));
  OR       g0784(.a(i_2_1_70_0), .b(i_2_1_46_0), .O(new_n801_));
  NOT      g0785(.a(new_n801_), .O(new_n802_));
  OR       g0786(.a(new_n802_), .b(new_n237_), .O(new_n803_));
  AND      g0787(.a(new_n803_), .b(new_n63_), .O(new_n804_));
  OR       g0788(.a(new_n804_), .b(new_n800_), .O(new_n805_));
  OR       g0789(.a(new_n805_), .b(new_n799_), .O(new_n806_));
  OR       g0790(.a(new_n806_), .b(new_n796_), .O(new_n807_));
  AND      g0791(.a(new_n807_), .b(i_2_1_13_0), .O(new_n808_));
  OR       g0792(.a(new_n808_), .b(new_n793_), .O(new_n809_));
  OR       g0793(.a(new_n809_), .b(new_n787_), .O(new_n810_));
  AND      g0794(.a(new_n810_), .b(i_2_1_38_0), .O(new_n811_));
  AND      g0795(.a(new_n644_), .b(i_2_1_68_0), .O(new_n812_));
  AND      g0796(.a(new_n636_), .b(new_n123_), .O(new_n813_));
  OR       g0797(.a(new_n813_), .b(new_n812_), .O(new_n814_));
  AND      g0798(.a(new_n814_), .b(i_2_1_41_0), .O(new_n815_));
  AND      g0799(.a(new_n575_), .b(i_2_1_70_0), .O(new_n816_));
  OR       g0800(.a(new_n816_), .b(new_n815_), .O(new_n817_));
  AND      g0801(.a(new_n817_), .b(new_n96_), .O(new_n818_));
  AND      g0802(.a(new_n127_), .b(new_n63_), .O(new_n819_));
  AND      g0803(.a(new_n819_), .b(new_n644_), .O(new_n820_));
  OR       g0804(.a(new_n84_), .b(new_n63_), .O(new_n821_));
  AND      g0805(.a(new_n821_), .b(new_n380_), .O(new_n822_));
  OR       g0806(.a(new_n822_), .b(new_n820_), .O(new_n823_));
  AND      g0807(.a(new_n823_), .b(i_2_1_68_0), .O(new_n824_));
  OR       g0808(.a(new_n489_), .b(new_n63_), .O(new_n825_));
  AND      g0809(.a(new_n825_), .b(new_n261_), .O(new_n826_));
  OR       g0810(.a(new_n691_), .b(new_n123_), .O(new_n827_));
  NAND     g0811(.a(new_n574_), .b(new_n28_), .O(new_n828_));
  AND      g0812(.a(new_n828_), .b(new_n636_), .O(new_n829_));
  AND      g0813(.a(new_n829_), .b(new_n827_), .O(new_n830_));
  OR       g0814(.a(new_n830_), .b(new_n826_), .O(new_n831_));
  OR       g0815(.a(new_n831_), .b(new_n824_), .O(new_n832_));
  OR       g0816(.a(new_n832_), .b(new_n818_), .O(new_n833_));
  AND      g0817(.a(new_n833_), .b(i_2_1_34_0), .O(new_n834_));
  NAND     g0818(.a(new_n574_), .b(new_n220_), .O(new_n835_));
  AND      g0819(.a(new_n835_), .b(i_2_1_13_0), .O(new_n836_));
  OR       g0820(.a(i_2_1_136_0), .b(i_2_1_41_0), .O(new_n837_));
  AND      g0821(.a(new_n338_), .b(i_2_1_68_0), .O(new_n838_));
  AND      g0822(.a(new_n838_), .b(new_n837_), .O(new_n839_));
  OR       g0823(.a(new_n839_), .b(new_n836_), .O(new_n840_));
  AND      g0824(.a(new_n840_), .b(i_2_1_135_0), .O(new_n841_));
  NAND     g0825(.a(new_n164_), .b(new_n28_), .O(new_n842_));
  OR       g0826(.a(new_n842_), .b(new_n838_), .O(new_n843_));
  AND      g0827(.a(new_n843_), .b(i_2_1_13_0), .O(new_n844_));
  OR       g0828(.a(new_n844_), .b(new_n841_), .O(new_n845_));
  AND      g0829(.a(new_n845_), .b(i_2_1_70_0), .O(new_n846_));
  AND      g0830(.a(new_n644_), .b(i_2_1_135_0), .O(new_n847_));
  NAND     g0831(.a(new_n847_), .b(new_n192_), .O(new_n848_));
  NAND     g0832(.a(new_n848_), .b(new_n625_), .O(new_n849_));
  AND      g0833(.a(new_n849_), .b(new_n431_), .O(new_n850_));
  OR       g0834(.a(new_n850_), .b(new_n846_), .O(new_n851_));
  OR       g0835(.a(new_n851_), .b(new_n834_), .O(new_n852_));
  OR       g0836(.a(new_n852_), .b(new_n811_), .O(new_n853_));
  OR       g0837(.a(new_n853_), .b(new_n759_), .O(new_n854_));
  OR       g0838(.a(new_n854_), .b(new_n683_), .O(new_n855_));
  AND      g0839(.a(new_n855_), .b(new_n32_), .O(new_n856_));
  OR       g0840(.a(new_n342_), .b(i_2_1_13_0), .O(new_n857_));
  OR       g0841(.a(new_n857_), .b(new_n797_), .O(new_n858_));
  AND      g0842(.a(new_n858_), .b(new_n798_), .O(new_n859_));
  OR       g0843(.a(new_n588_), .b(i_2_1_34_0), .O(new_n860_));
  OR       g0844(.a(i_2_1_70_0), .b(i_2_1_41_0), .O(new_n861_));
  NOT      g0845(.a(new_n861_), .O(new_n862_));
  AND      g0846(.a(new_n862_), .b(new_n860_), .O(new_n863_));
  OR       g0847(.a(new_n863_), .b(new_n859_), .O(new_n864_));
  AND      g0848(.a(new_n864_), .b(i_2_1_32_0), .O(new_n865_));
  OR       g0849(.a(new_n697_), .b(i_2_1_41_0), .O(new_n866_));
  AND      g0850(.a(new_n866_), .b(new_n575_), .O(new_n867_));
  OR       g0851(.a(new_n438_), .b(new_n237_), .O(new_n868_));
  AND      g0852(.a(new_n868_), .b(new_n63_), .O(new_n869_));
  OR       g0853(.a(new_n567_), .b(new_n397_), .O(new_n870_));
  AND      g0854(.a(new_n870_), .b(new_n272_), .O(new_n871_));
  OR       g0855(.a(new_n871_), .b(new_n869_), .O(new_n872_));
  OR       g0856(.a(new_n872_), .b(new_n867_), .O(new_n873_));
  OR       g0857(.a(new_n873_), .b(new_n865_), .O(new_n874_));
  AND      g0858(.a(new_n874_), .b(i_2_1_135_0), .O(new_n875_));
  OR       g0859(.a(new_n397_), .b(new_n141_), .O(new_n876_));
  AND      g0860(.a(new_n876_), .b(i_2_1_68_0), .O(new_n877_));
  OR       g0861(.a(new_n337_), .b(new_n32_), .O(new_n878_));
  NAND     g0862(.a(new_n594_), .b(i_2_1_13_0), .O(new_n879_));
  AND      g0863(.a(new_n879_), .b(new_n34_), .O(new_n880_));
  NAND     g0864(.a(new_n880_), .b(new_n878_), .O(new_n881_));
  AND      g0865(.a(new_n881_), .b(new_n54_), .O(new_n882_));
  OR       g0866(.a(new_n882_), .b(new_n877_), .O(new_n883_));
  AND      g0867(.a(new_n883_), .b(i_2_1_41_0), .O(new_n884_));
  OR       g0868(.a(new_n19_), .b(i_2_1_32_0), .O(new_n885_));
  AND      g0869(.a(new_n885_), .b(i_2_1_13_0), .O(new_n886_));
  AND      g0870(.a(new_n802_), .b(i_2_1_32_0), .O(new_n887_));
  OR       g0871(.a(new_n887_), .b(new_n886_), .O(new_n888_));
  AND      g0872(.a(new_n888_), .b(new_n63_), .O(new_n889_));
  AND      g0873(.a(new_n798_), .b(i_2_1_32_0), .O(new_n890_));
  NOT      g0874(.a(new_n838_), .O(new_n891_));
  NOT      g0875(.a(i_2_1_32_0), .O(new_n892_));
  AND      g0876(.a(i_2_1_49_0), .b(new_n892_), .O(new_n893_));
  OR       g0877(.a(new_n893_), .b(new_n531_), .O(new_n894_));
  NAND     g0878(.a(new_n894_), .b(new_n891_), .O(new_n895_));
  OR       g0879(.a(new_n895_), .b(new_n890_), .O(new_n896_));
  AND      g0880(.a(new_n896_), .b(i_2_1_70_0), .O(new_n897_));
  OR       g0881(.a(new_n897_), .b(new_n889_), .O(new_n898_));
  OR       g0882(.a(new_n898_), .b(new_n884_), .O(new_n899_));
  OR       g0883(.a(new_n899_), .b(new_n875_), .O(new_n900_));
  AND      g0884(.a(new_n900_), .b(i_2_1_136_0), .O(new_n901_));
  OR       g0885(.a(new_n397_), .b(new_n347_), .O(new_n902_));
  AND      g0886(.a(new_n19_), .b(i_2_1_32_0), .O(new_n903_));
  OR       g0887(.a(new_n489_), .b(i_2_1_41_0), .O(new_n904_));
  OR       g0888(.a(new_n904_), .b(new_n903_), .O(new_n905_));
  AND      g0889(.a(new_n905_), .b(new_n902_), .O(new_n906_));
  OR       g0890(.a(new_n906_), .b(new_n645_), .O(new_n907_));
  AND      g0891(.a(new_n907_), .b(i_2_1_68_0), .O(new_n908_));
  AND      g0892(.a(new_n403_), .b(i_2_1_13_0), .O(new_n909_));
  AND      g0893(.a(i_2_1_70_0), .b(i_2_1_32_0), .O(new_n910_));
  AND      g0894(.a(new_n910_), .b(i_2_1_54_0), .O(new_n911_));
  OR       g0895(.a(new_n911_), .b(new_n535_), .O(new_n912_));
  OR       g0896(.a(new_n912_), .b(new_n909_), .O(new_n913_));
  OR       g0897(.a(i_2_1_136_0), .b(new_n32_), .O(new_n914_));
  OR       g0898(.a(new_n446_), .b(i_2_1_46_0), .O(new_n915_));
  OR       g0899(.a(new_n915_), .b(new_n914_), .O(new_n916_));
  NAND     g0900(.a(new_n916_), .b(new_n57_), .O(new_n917_));
  OR       g0901(.a(new_n917_), .b(new_n913_), .O(new_n918_));
  AND      g0902(.a(new_n918_), .b(i_2_1_41_0), .O(new_n919_));
  OR       g0903(.a(new_n261_), .b(i_2_1_135_0), .O(new_n920_));
  OR       g0904(.a(new_n123_), .b(i_2_1_32_0), .O(new_n921_));
  OR       g0905(.a(new_n802_), .b(new_n272_), .O(new_n922_));
  AND      g0906(.a(new_n922_), .b(new_n921_), .O(new_n923_));
  AND      g0907(.a(new_n923_), .b(new_n920_), .O(new_n924_));
  OR       g0908(.a(new_n924_), .b(new_n919_), .O(new_n925_));
  OR       g0909(.a(new_n925_), .b(new_n908_), .O(new_n926_));
  AND      g0910(.a(new_n926_), .b(new_n63_), .O(new_n927_));
  AND      g0911(.a(new_n176_), .b(i_2_1_32_0), .O(new_n928_));
  OR       g0912(.a(new_n928_), .b(new_n470_), .O(new_n929_));
  AND      g0913(.a(new_n885_), .b(new_n237_), .O(new_n930_));
  OR       g0914(.a(new_n930_), .b(new_n835_), .O(new_n931_));
  AND      g0915(.a(new_n931_), .b(new_n929_), .O(new_n932_));
  AND      g0916(.a(new_n27_), .b(i_2_1_34_0), .O(new_n933_));
  OR       g0917(.a(new_n933_), .b(new_n445_), .O(new_n934_));
  AND      g0918(.a(new_n934_), .b(i_2_1_32_0), .O(new_n935_));
  NOT      g0919(.a(new_n96_), .O(new_n936_));
  AND      g0920(.a(new_n567_), .b(new_n936_), .O(new_n937_));
  OR       g0921(.a(new_n937_), .b(new_n935_), .O(new_n938_));
  AND      g0922(.a(new_n938_), .b(i_2_1_135_0), .O(new_n939_));
  NAND     g0923(.a(new_n574_), .b(new_n52_), .O(new_n940_));
  AND      g0924(.a(new_n940_), .b(i_2_1_13_0), .O(new_n941_));
  OR       g0925(.a(new_n941_), .b(new_n930_), .O(new_n942_));
  OR       g0926(.a(new_n942_), .b(new_n939_), .O(new_n943_));
  AND      g0927(.a(new_n943_), .b(i_2_1_70_0), .O(new_n944_));
  OR       g0928(.a(new_n944_), .b(new_n932_), .O(new_n945_));
  OR       g0929(.a(new_n945_), .b(new_n927_), .O(new_n946_));
  OR       g0930(.a(new_n946_), .b(new_n901_), .O(new_n947_));
  AND      g0931(.a(new_n947_), .b(new_n20_), .O(new_n948_));
  OR       g0932(.a(new_n762_), .b(i_2_1_135_0), .O(new_n949_));
  AND      g0933(.a(new_n949_), .b(new_n19_), .O(new_n950_));
  NAND     g0934(.a(new_n94_), .b(new_n220_), .O(new_n951_));
  AND      g0935(.a(new_n951_), .b(i_2_1_32_0), .O(new_n952_));
  AND      g0936(.a(i_2_1_136_0), .b(i_2_1_57_0), .O(new_n953_));
  NOT      g0937(.a(new_n953_), .O(new_n954_));
  OR       g0938(.a(new_n954_), .b(new_n762_), .O(new_n955_));
  NAND     g0939(.a(new_n955_), .b(new_n879_), .O(new_n956_));
  OR       g0940(.a(new_n956_), .b(new_n952_), .O(new_n957_));
  OR       g0941(.a(new_n957_), .b(new_n950_), .O(new_n958_));
  AND      g0942(.a(new_n958_), .b(i_2_1_34_0), .O(new_n959_));
  OR       g0943(.a(new_n364_), .b(new_n19_), .O(new_n960_));
  AND      g0944(.a(new_n960_), .b(new_n63_), .O(new_n961_));
  OR       g0945(.a(new_n445_), .b(new_n21_), .O(new_n962_));
  OR       g0946(.a(new_n19_), .b(i_2_1_41_0), .O(new_n963_));
  AND      g0947(.a(new_n963_), .b(i_2_1_136_0), .O(new_n964_));
  OR       g0948(.a(new_n964_), .b(new_n962_), .O(new_n965_));
  OR       g0949(.a(new_n965_), .b(new_n961_), .O(new_n966_));
  AND      g0950(.a(new_n966_), .b(i_2_1_13_0), .O(new_n967_));
  AND      g0951(.a(new_n127_), .b(new_n19_), .O(new_n968_));
  AND      g0952(.a(new_n968_), .b(new_n321_), .O(new_n969_));
  OR       g0953(.a(new_n760_), .b(new_n63_), .O(new_n970_));
  AND      g0954(.a(new_n970_), .b(new_n969_), .O(new_n971_));
  OR       g0955(.a(new_n380_), .b(new_n148_), .O(new_n972_));
  AND      g0956(.a(new_n972_), .b(i_2_1_32_0), .O(new_n973_));
  OR       g0957(.a(new_n973_), .b(new_n971_), .O(new_n974_));
  OR       g0958(.a(new_n974_), .b(new_n967_), .O(new_n975_));
  OR       g0959(.a(new_n975_), .b(new_n959_), .O(new_n976_));
  AND      g0960(.a(new_n976_), .b(i_2_1_70_0), .O(new_n977_));
  OR       g0961(.a(new_n337_), .b(new_n54_), .O(new_n978_));
  NAND     g0962(.a(new_n978_), .b(new_n780_), .O(new_n979_));
  AND      g0963(.a(new_n979_), .b(i_2_1_32_0), .O(new_n980_));
  AND      g0964(.a(new_n489_), .b(new_n365_), .O(new_n981_));
  OR       g0965(.a(new_n595_), .b(new_n380_), .O(new_n982_));
  OR       g0966(.a(new_n364_), .b(i_2_1_32_0), .O(new_n983_));
  AND      g0967(.a(new_n983_), .b(new_n982_), .O(new_n984_));
  OR       g0968(.a(new_n984_), .b(new_n981_), .O(new_n985_));
  OR       g0969(.a(new_n985_), .b(new_n980_), .O(new_n986_));
  AND      g0970(.a(new_n986_), .b(i_2_1_136_0), .O(new_n987_));
  OR       g0971(.a(i_2_1_41_0), .b(i_2_1_13_0), .O(new_n988_));
  AND      g0972(.a(new_n988_), .b(i_2_1_34_0), .O(new_n989_));
  OR       g0973(.a(new_n347_), .b(i_2_1_32_0), .O(new_n990_));
  OR       g0974(.a(new_n990_), .b(new_n989_), .O(new_n991_));
  AND      g0975(.a(new_n638_), .b(new_n338_), .O(new_n992_));
  AND      g0976(.a(new_n992_), .b(new_n991_), .O(new_n993_));
  AND      g0977(.a(i_2_1_57_0), .b(i_2_1_51_0), .O(new_n994_));
  OR       g0978(.a(new_n994_), .b(new_n21_), .O(new_n995_));
  AND      g0979(.a(new_n995_), .b(i_2_1_32_0), .O(new_n996_));
  AND      g0980(.a(new_n996_), .b(new_n800_), .O(new_n997_));
  OR       g0981(.a(new_n997_), .b(new_n993_), .O(new_n998_));
  OR       g0982(.a(new_n998_), .b(new_n987_), .O(new_n999_));
  OR       g0983(.a(new_n999_), .b(new_n977_), .O(new_n1000_));
  AND      g0984(.a(new_n1000_), .b(i_2_1_68_0), .O(new_n1001_));
  NAND     g0985(.a(new_n438_), .b(new_n54_), .O(new_n1002_));
  NAND     g0986(.a(new_n1002_), .b(new_n481_), .O(new_n1003_));
  AND      g0987(.a(new_n1003_), .b(i_2_1_136_0), .O(new_n1004_));
  AND      g0988(.a(new_n123_), .b(new_n27_), .O(new_n1005_));
  AND      g0989(.a(new_n1005_), .b(i_2_1_41_0), .O(new_n1006_));
  OR       g0990(.a(new_n953_), .b(i_2_1_13_0), .O(new_n1007_));
  AND      g0991(.a(new_n1007_), .b(i_2_1_32_0), .O(new_n1008_));
  OR       g0992(.a(new_n1008_), .b(new_n1006_), .O(new_n1009_));
  OR       g0993(.a(new_n1009_), .b(new_n1004_), .O(new_n1010_));
  AND      g0994(.a(new_n1010_), .b(new_n63_), .O(new_n1011_));
  OR       g0995(.a(new_n1011_), .b(new_n388_), .O(new_n1012_));
  AND      g0996(.a(new_n1012_), .b(i_2_1_34_0), .O(new_n1013_));
  AND      g0997(.a(new_n996_), .b(new_n794_), .O(new_n1014_));
  AND      g0998(.a(new_n446_), .b(new_n63_), .O(new_n1015_));
  NAND     g0999(.a(new_n1015_), .b(new_n712_), .O(new_n1016_));
  AND      g1000(.a(new_n53_), .b(i_2_1_34_0), .O(new_n1017_));
  NAND     g1001(.a(new_n1017_), .b(i_2_1_57_0), .O(new_n1018_));
  OR       g1002(.a(new_n1018_), .b(new_n54_), .O(new_n1019_));
  NAND     g1003(.a(new_n1019_), .b(new_n1016_), .O(new_n1020_));
  OR       g1004(.a(new_n1020_), .b(new_n1014_), .O(new_n1021_));
  AND      g1005(.a(new_n1021_), .b(i_2_1_13_0), .O(new_n1022_));
  AND      g1006(.a(new_n606_), .b(i_2_1_135_0), .O(new_n1023_));
  NOT      g1007(.a(new_n51_), .O(new_n1024_));
  AND      g1008(.a(new_n1024_), .b(i_2_1_32_0), .O(new_n1025_));
  AND      g1009(.a(new_n1025_), .b(new_n165_), .O(new_n1026_));
  AND      g1010(.a(new_n124_), .b(i_2_1_34_0), .O(new_n1027_));
  OR       g1011(.a(new_n1027_), .b(new_n1026_), .O(new_n1028_));
  AND      g1012(.a(new_n1028_), .b(i_2_1_41_0), .O(new_n1029_));
  OR       g1013(.a(new_n1029_), .b(new_n1023_), .O(new_n1030_));
  OR       g1014(.a(new_n1030_), .b(new_n1022_), .O(new_n1031_));
  AND      g1015(.a(new_n1031_), .b(new_n19_), .O(new_n1032_));
  AND      g1016(.a(new_n362_), .b(i_2_1_13_0), .O(new_n1033_));
  OR       g1017(.a(new_n1033_), .b(new_n309_), .O(new_n1034_));
  AND      g1018(.a(new_n1034_), .b(new_n910_), .O(new_n1035_));
  OR       g1019(.a(new_n1035_), .b(new_n1032_), .O(new_n1036_));
  OR       g1020(.a(new_n1036_), .b(new_n1013_), .O(new_n1037_));
  OR       g1021(.a(new_n1037_), .b(new_n1001_), .O(new_n1038_));
  OR       g1022(.a(new_n1038_), .b(new_n948_), .O(new_n1039_));
  AND      g1023(.a(new_n1039_), .b(i_2_1_38_0), .O(new_n1040_));
  OR       g1024(.a(new_n103_), .b(i_2_1_57_0), .O(new_n1041_));
  NAND     g1025(.a(new_n399_), .b(i_2_1_46_0), .O(new_n1042_));
  AND      g1026(.a(new_n1042_), .b(i_2_1_41_0), .O(new_n1043_));
  AND      g1027(.a(new_n1043_), .b(new_n1041_), .O(new_n1044_));
  AND      g1028(.a(new_n257_), .b(i_2_1_34_0), .O(new_n1045_));
  AND      g1029(.a(new_n575_), .b(new_n65_), .O(new_n1046_));
  AND      g1030(.a(new_n636_), .b(i_2_1_70_0), .O(new_n1047_));
  OR       g1031(.a(new_n1047_), .b(new_n1046_), .O(new_n1048_));
  OR       g1032(.a(new_n1048_), .b(new_n1045_), .O(new_n1049_));
  OR       g1033(.a(new_n1049_), .b(new_n1044_), .O(new_n1050_));
  AND      g1034(.a(new_n1050_), .b(new_n63_), .O(new_n1051_));
  NOT      g1035(.a(new_n436_), .O(new_n1052_));
  OR       g1036(.a(new_n720_), .b(new_n1052_), .O(new_n1053_));
  AND      g1037(.a(new_n1053_), .b(i_2_1_135_0), .O(new_n1054_));
  NAND     g1038(.a(new_n436_), .b(new_n53_), .O(new_n1055_));
  AND      g1039(.a(new_n1055_), .b(i_2_1_41_0), .O(new_n1056_));
  OR       g1040(.a(new_n1056_), .b(new_n1054_), .O(new_n1057_));
  AND      g1041(.a(new_n1057_), .b(i_2_1_68_0), .O(new_n1058_));
  OR       g1042(.a(new_n438_), .b(i_2_1_57_0), .O(new_n1059_));
  AND      g1043(.a(new_n868_), .b(i_2_1_49_0), .O(new_n1060_));
  AND      g1044(.a(new_n1060_), .b(new_n1059_), .O(new_n1061_));
  OR       g1045(.a(new_n1061_), .b(new_n1058_), .O(new_n1062_));
  OR       g1046(.a(new_n1062_), .b(new_n1051_), .O(new_n1063_));
  AND      g1047(.a(new_n1063_), .b(i_2_1_136_0), .O(new_n1064_));
  NOT      g1048(.a(new_n399_), .O(new_n1065_));
  AND      g1049(.a(new_n838_), .b(new_n1065_), .O(new_n1066_));
  AND      g1050(.a(new_n684_), .b(new_n20_), .O(new_n1067_));
  NOT      g1051(.a(new_n169_), .O(new_n1068_));
  AND      g1052(.a(new_n575_), .b(new_n1068_), .O(new_n1069_));
  OR       g1053(.a(new_n1069_), .b(new_n1067_), .O(new_n1070_));
  OR       g1054(.a(i_2_1_68_0), .b(new_n220_), .O(new_n1071_));
  NAND     g1055(.a(new_n1071_), .b(new_n53_), .O(new_n1072_));
  AND      g1056(.a(new_n1072_), .b(new_n63_), .O(new_n1073_));
  NAND     g1057(.a(i_2_1_51_0), .b(i_2_1_49_0), .O(new_n1074_));
  NOT      g1058(.a(new_n1074_), .O(new_n1075_));
  OR       g1059(.a(new_n1075_), .b(new_n175_), .O(new_n1076_));
  AND      g1060(.a(new_n1076_), .b(i_2_1_41_0), .O(new_n1077_));
  OR       g1061(.a(new_n1077_), .b(new_n1073_), .O(new_n1078_));
  OR       g1062(.a(new_n1078_), .b(new_n1070_), .O(new_n1079_));
  AND      g1063(.a(new_n1079_), .b(i_2_1_34_0), .O(new_n1080_));
  OR       g1064(.a(new_n1080_), .b(new_n1066_), .O(new_n1081_));
  OR       g1065(.a(new_n1081_), .b(new_n1064_), .O(new_n1082_));
  AND      g1066(.a(new_n1082_), .b(i_2_1_32_0), .O(new_n1083_));
  AND      g1067(.a(new_n575_), .b(new_n96_), .O(new_n1084_));
  OR       g1068(.a(new_n141_), .b(new_n20_), .O(new_n1085_));
  AND      g1069(.a(new_n1085_), .b(new_n27_), .O(new_n1086_));
  OR       g1070(.a(new_n1086_), .b(new_n1084_), .O(new_n1087_));
  AND      g1071(.a(new_n1087_), .b(i_2_1_135_0), .O(new_n1088_));
  NAND     g1072(.a(new_n574_), .b(i_2_1_57_0), .O(new_n1089_));
  AND      g1073(.a(new_n1089_), .b(new_n607_), .O(new_n1090_));
  OR       g1074(.a(new_n1090_), .b(new_n243_), .O(new_n1091_));
  OR       g1075(.a(new_n1091_), .b(new_n1088_), .O(new_n1092_));
  AND      g1076(.a(new_n1092_), .b(i_2_1_41_0), .O(new_n1093_));
  AND      g1077(.a(new_n362_), .b(new_n338_), .O(new_n1094_));
  OR       g1078(.a(new_n1052_), .b(new_n364_), .O(new_n1095_));
  OR       g1079(.a(new_n1095_), .b(new_n1094_), .O(new_n1096_));
  AND      g1080(.a(new_n1096_), .b(i_2_1_68_0), .O(new_n1097_));
  OR       g1081(.a(new_n1097_), .b(new_n1067_), .O(new_n1098_));
  AND      g1082(.a(new_n1098_), .b(i_2_1_32_0), .O(new_n1099_));
  AND      g1083(.a(new_n74_), .b(i_2_1_136_0), .O(new_n1100_));
  AND      g1084(.a(new_n127_), .b(i_2_1_34_0), .O(new_n1101_));
  OR       g1085(.a(new_n1101_), .b(new_n63_), .O(new_n1102_));
  AND      g1086(.a(new_n794_), .b(new_n19_), .O(new_n1103_));
  AND      g1087(.a(new_n1103_), .b(new_n1102_), .O(new_n1104_));
  OR       g1088(.a(new_n1104_), .b(new_n1100_), .O(new_n1105_));
  AND      g1089(.a(new_n1105_), .b(i_2_1_68_0), .O(new_n1106_));
  NAND     g1090(.a(new_n237_), .b(i_2_1_49_0), .O(new_n1107_));
  OR       g1091(.a(new_n337_), .b(new_n164_), .O(new_n1108_));
  NAND     g1092(.a(new_n1108_), .b(new_n1107_), .O(new_n1109_));
  AND      g1093(.a(new_n1109_), .b(new_n20_), .O(new_n1110_));
  OR       g1094(.a(new_n1110_), .b(new_n1106_), .O(new_n1111_));
  OR       g1095(.a(new_n1111_), .b(new_n1099_), .O(new_n1112_));
  OR       g1096(.a(new_n1112_), .b(new_n1093_), .O(new_n1113_));
  AND      g1097(.a(new_n1113_), .b(i_2_1_70_0), .O(new_n1114_));
  AND      g1098(.a(new_n797_), .b(new_n191_), .O(new_n1115_));
  OR       g1099(.a(new_n669_), .b(new_n20_), .O(new_n1116_));
  AND      g1100(.a(new_n1116_), .b(i_2_1_41_0), .O(new_n1117_));
  OR       g1101(.a(new_n28_), .b(i_2_1_46_0), .O(new_n1118_));
  NAND     g1102(.a(new_n1118_), .b(i_2_1_57_0), .O(new_n1119_));
  AND      g1103(.a(new_n1119_), .b(new_n828_), .O(new_n1120_));
  OR       g1104(.a(new_n1120_), .b(new_n1117_), .O(new_n1121_));
  AND      g1105(.a(new_n1121_), .b(i_2_1_34_0), .O(new_n1122_));
  AND      g1106(.a(new_n762_), .b(i_2_1_136_0), .O(new_n1123_));
  AND      g1107(.a(new_n1123_), .b(new_n257_), .O(new_n1124_));
  AND      g1108(.a(new_n1124_), .b(new_n1069_), .O(new_n1125_));
  OR       g1109(.a(new_n1125_), .b(new_n1122_), .O(new_n1126_));
  AND      g1110(.a(new_n1126_), .b(i_2_1_135_0), .O(new_n1127_));
  OR       g1111(.a(new_n1127_), .b(new_n1115_), .O(new_n1128_));
  OR       g1112(.a(new_n1128_), .b(new_n1114_), .O(new_n1129_));
  OR       g1113(.a(new_n1129_), .b(new_n1083_), .O(new_n1130_));
  AND      g1114(.a(new_n1130_), .b(i_2_1_13_0), .O(new_n1131_));
  OR       g1115(.a(i_2_1_135_0), .b(new_n18_), .O(new_n1132_));
  NAND     g1116(.a(new_n1132_), .b(new_n26_), .O(new_n1133_));
  AND      g1117(.a(new_n1133_), .b(i_2_1_32_0), .O(new_n1134_));
  OR       g1118(.a(new_n1134_), .b(new_n397_), .O(new_n1135_));
  AND      g1119(.a(new_n1135_), .b(new_n20_), .O(new_n1136_));
  AND      g1120(.a(new_n84_), .b(i_2_1_68_0), .O(new_n1137_));
  OR       g1121(.a(new_n123_), .b(new_n63_), .O(new_n1138_));
  AND      g1122(.a(new_n1138_), .b(new_n1137_), .O(new_n1139_));
  OR       g1123(.a(new_n1132_), .b(new_n53_), .O(new_n1140_));
  NAND     g1124(.a(new_n1140_), .b(i_2_1_49_0), .O(new_n1141_));
  AND      g1125(.a(new_n1141_), .b(i_2_1_32_0), .O(new_n1142_));
  OR       g1126(.a(new_n1142_), .b(new_n1139_), .O(new_n1143_));
  AND      g1127(.a(new_n1143_), .b(new_n19_), .O(new_n1144_));
  OR       g1128(.a(new_n1144_), .b(new_n1136_), .O(new_n1145_));
  AND      g1129(.a(new_n1145_), .b(i_2_1_136_0), .O(new_n1146_));
  AND      g1130(.a(new_n1089_), .b(i_2_1_32_0), .O(new_n1147_));
  OR       g1131(.a(new_n838_), .b(new_n194_), .O(new_n1148_));
  AND      g1132(.a(new_n1148_), .b(i_2_1_135_0), .O(new_n1149_));
  OR       g1133(.a(new_n1149_), .b(new_n1147_), .O(new_n1150_));
  AND      g1134(.a(new_n1150_), .b(i_2_1_70_0), .O(new_n1151_));
  AND      g1135(.a(new_n414_), .b(new_n77_), .O(new_n1152_));
  AND      g1136(.a(new_n1152_), .b(new_n893_), .O(new_n1153_));
  OR       g1137(.a(new_n1153_), .b(new_n1151_), .O(new_n1154_));
  OR       g1138(.a(new_n1154_), .b(new_n1146_), .O(new_n1155_));
  AND      g1139(.a(new_n1155_), .b(i_2_1_41_0), .O(new_n1156_));
  AND      g1140(.a(i_2_1_135_0), .b(i_2_1_32_0), .O(new_n1157_));
  NOT      g1141(.a(new_n1157_), .O(new_n1158_));
  OR       g1142(.a(new_n337_), .b(i_2_1_57_0), .O(new_n1159_));
  OR       g1143(.a(new_n1159_), .b(new_n1158_), .O(new_n1160_));
  OR       g1144(.a(new_n903_), .b(i_2_1_136_0), .O(new_n1161_));
  AND      g1145(.a(new_n1161_), .b(new_n20_), .O(new_n1162_));
  OR       g1146(.a(new_n20_), .b(i_2_1_32_0), .O(new_n1163_));
  AND      g1147(.a(new_n1163_), .b(new_n493_), .O(new_n1164_));
  AND      g1148(.a(new_n489_), .b(i_2_1_136_0), .O(new_n1165_));
  AND      g1149(.a(i_2_1_136_0), .b(i_2_1_32_0), .O(new_n1166_));
  OR       g1150(.a(new_n1166_), .b(new_n1165_), .O(new_n1167_));
  OR       g1151(.a(new_n1167_), .b(new_n1164_), .O(new_n1168_));
  AND      g1152(.a(new_n1168_), .b(i_2_1_68_0), .O(new_n1169_));
  OR       g1153(.a(new_n1169_), .b(new_n1162_), .O(new_n1170_));
  AND      g1154(.a(new_n1170_), .b(new_n63_), .O(new_n1171_));
  AND      g1155(.a(new_n131_), .b(i_2_1_32_0), .O(new_n1172_));
  OR       g1156(.a(new_n1172_), .b(new_n1171_), .O(new_n1173_));
  NAND     g1157(.a(new_n1173_), .b(i_2_1_70_0), .O(new_n1174_));
  NAND     g1158(.a(new_n1174_), .b(new_n1160_), .O(new_n1175_));
  OR       g1159(.a(new_n1175_), .b(new_n1156_), .O(new_n1176_));
  AND      g1160(.a(new_n1176_), .b(i_2_1_34_0), .O(new_n1177_));
  AND      g1161(.a(new_n438_), .b(new_n65_), .O(new_n1178_));
  OR       g1162(.a(new_n760_), .b(new_n353_), .O(new_n1179_));
  AND      g1163(.a(new_n1179_), .b(new_n20_), .O(new_n1180_));
  OR       g1164(.a(new_n1180_), .b(new_n1178_), .O(new_n1181_));
  AND      g1165(.a(new_n1181_), .b(new_n63_), .O(new_n1182_));
  AND      g1166(.a(new_n257_), .b(new_n124_), .O(new_n1183_));
  OR       g1167(.a(new_n1183_), .b(new_n1182_), .O(new_n1184_));
  AND      g1168(.a(new_n1184_), .b(i_2_1_32_0), .O(new_n1185_));
  AND      g1169(.a(new_n342_), .b(new_n129_), .O(new_n1186_));
  OR       g1170(.a(new_n1186_), .b(new_n1185_), .O(new_n1187_));
  AND      g1171(.a(new_n1187_), .b(new_n575_), .O(new_n1188_));
  OR       g1172(.a(new_n39_), .b(new_n19_), .O(new_n1189_));
  AND      g1173(.a(new_n1157_), .b(new_n438_), .O(new_n1190_));
  AND      g1174(.a(new_n1190_), .b(new_n190_), .O(new_n1191_));
  AND      g1175(.a(new_n1191_), .b(new_n1189_), .O(new_n1192_));
  OR       g1176(.a(new_n1192_), .b(new_n1188_), .O(new_n1193_));
  OR       g1177(.a(new_n1193_), .b(new_n1177_), .O(new_n1194_));
  OR       g1178(.a(new_n1194_), .b(new_n1131_), .O(new_n1195_));
  OR       g1179(.a(new_n1195_), .b(new_n1040_), .O(new_n1196_));
  OR       g1180(.a(new_n1196_), .b(new_n856_), .O(new_n1197_));
  OR       g1181(.a(new_n1197_), .b(new_n562_), .O(new_n1198_));
  AND      g1182(.a(new_n1198_), .b(new_n17_), .O(new_n1199_));
  AND      g1183(.a(new_n580_), .b(i_2_1_34_0), .O(new_n1200_));
  OR       g1184(.a(new_n362_), .b(new_n73_), .O(new_n1201_));
  AND      g1185(.a(new_n1201_), .b(new_n19_), .O(new_n1202_));
  OR       g1186(.a(new_n1202_), .b(new_n1200_), .O(new_n1203_));
  AND      g1187(.a(new_n1203_), .b(i_2_1_136_0), .O(new_n1204_));
  NAND     g1188(.a(new_n37_), .b(new_n27_), .O(new_n1205_));
  NAND     g1189(.a(new_n1205_), .b(new_n704_), .O(new_n1206_));
  AND      g1190(.a(new_n1206_), .b(new_n220_), .O(new_n1207_));
  OR       g1191(.a(new_n431_), .b(i_2_1_34_0), .O(new_n1208_));
  AND      g1192(.a(new_n54_), .b(i_2_1_70_0), .O(new_n1209_));
  AND      g1193(.a(new_n283_), .b(i_2_1_68_0), .O(new_n1210_));
  OR       g1194(.a(new_n1210_), .b(new_n1209_), .O(new_n1211_));
  AND      g1195(.a(new_n1211_), .b(new_n1208_), .O(new_n1212_));
  AND      g1196(.a(new_n74_), .b(i_2_1_41_0), .O(new_n1213_));
  OR       g1197(.a(i_2_1_38_0), .b(i_2_1_34_0), .O(new_n1214_));
  OR       g1198(.a(new_n1214_), .b(i_2_1_41_0), .O(new_n1215_));
  AND      g1199(.a(new_n1215_), .b(new_n176_), .O(new_n1216_));
  OR       g1200(.a(new_n1216_), .b(new_n1213_), .O(new_n1217_));
  OR       g1201(.a(new_n1217_), .b(new_n1212_), .O(new_n1218_));
  OR       g1202(.a(new_n1218_), .b(new_n1207_), .O(new_n1219_));
  OR       g1203(.a(new_n1219_), .b(new_n1204_), .O(new_n1220_));
  AND      g1204(.a(new_n1220_), .b(new_n18_), .O(new_n1221_));
  OR       g1205(.a(new_n569_), .b(new_n265_), .O(new_n1222_));
  OR       g1206(.a(new_n364_), .b(i_2_1_68_0), .O(new_n1223_));
  AND      g1207(.a(new_n1223_), .b(i_2_1_38_0), .O(new_n1224_));
  AND      g1208(.a(new_n1224_), .b(new_n1222_), .O(new_n1225_));
  AND      g1209(.a(new_n870_), .b(i_2_1_70_0), .O(new_n1226_));
  OR       g1210(.a(new_n1226_), .b(new_n445_), .O(new_n1227_));
  AND      g1211(.a(new_n1227_), .b(i_2_1_135_0), .O(new_n1228_));
  OR       g1212(.a(new_n574_), .b(i_2_1_135_0), .O(new_n1229_));
  NAND     g1213(.a(new_n1229_), .b(new_n780_), .O(new_n1230_));
  AND      g1214(.a(new_n1230_), .b(i_2_1_51_0), .O(new_n1231_));
  OR       g1215(.a(new_n660_), .b(i_2_1_34_0), .O(new_n1232_));
  AND      g1216(.a(new_n1232_), .b(i_2_1_13_0), .O(new_n1233_));
  OR       g1217(.a(new_n1233_), .b(new_n1231_), .O(new_n1234_));
  OR       g1218(.a(new_n1234_), .b(new_n1228_), .O(new_n1235_));
  OR       g1219(.a(new_n1235_), .b(new_n1225_), .O(new_n1236_));
  AND      g1220(.a(new_n1236_), .b(i_2_1_136_0), .O(new_n1237_));
  OR       g1221(.a(new_n470_), .b(new_n273_), .O(new_n1238_));
  AND      g1222(.a(new_n1238_), .b(i_2_1_135_0), .O(new_n1239_));
  OR       g1223(.a(new_n532_), .b(new_n19_), .O(new_n1240_));
  OR       g1224(.a(new_n175_), .b(i_2_1_41_0), .O(new_n1241_));
  OR       g1225(.a(new_n644_), .b(i_2_1_34_0), .O(new_n1242_));
  AND      g1226(.a(new_n1242_), .b(new_n1241_), .O(new_n1243_));
  OR       g1227(.a(new_n1243_), .b(i_2_1_70_0), .O(new_n1244_));
  AND      g1228(.a(new_n1244_), .b(new_n1240_), .O(new_n1245_));
  OR       g1229(.a(new_n1245_), .b(new_n1239_), .O(new_n1246_));
  AND      g1230(.a(new_n1246_), .b(i_2_1_68_0), .O(new_n1247_));
  AND      g1231(.a(new_n387_), .b(i_2_1_34_0), .O(new_n1248_));
  OR       g1232(.a(new_n279_), .b(i_2_1_13_0), .O(new_n1249_));
  AND      g1233(.a(new_n1249_), .b(new_n963_), .O(new_n1250_));
  AND      g1234(.a(new_n74_), .b(i_2_1_51_0), .O(new_n1251_));
  OR       g1235(.a(new_n1251_), .b(new_n445_), .O(new_n1252_));
  OR       g1236(.a(new_n1252_), .b(new_n1250_), .O(new_n1253_));
  AND      g1237(.a(new_n1253_), .b(i_2_1_70_0), .O(new_n1254_));
  OR       g1238(.a(new_n1254_), .b(new_n1248_), .O(new_n1255_));
  OR       g1239(.a(new_n1255_), .b(new_n1247_), .O(new_n1256_));
  OR       g1240(.a(new_n1256_), .b(new_n1237_), .O(new_n1257_));
  OR       g1241(.a(new_n1257_), .b(new_n1221_), .O(new_n1258_));
  AND      g1242(.a(new_n1258_), .b(new_n20_), .O(new_n1259_));
  AND      g1243(.a(new_n1132_), .b(i_2_1_38_0), .O(new_n1260_));
  AND      g1244(.a(new_n362_), .b(new_n18_), .O(new_n1261_));
  OR       g1245(.a(new_n1261_), .b(new_n644_), .O(new_n1262_));
  OR       g1246(.a(new_n1262_), .b(new_n1260_), .O(new_n1263_));
  AND      g1247(.a(new_n1263_), .b(i_2_1_34_0), .O(new_n1264_));
  AND      g1248(.a(new_n18_), .b(i_2_1_41_0), .O(new_n1265_));
  AND      g1249(.a(new_n1265_), .b(i_2_1_136_0), .O(new_n1266_));
  NOT      g1250(.a(new_n287_), .O(new_n1267_));
  NOT      g1251(.a(new_n364_), .O(new_n1268_));
  OR       g1252(.a(new_n389_), .b(new_n1268_), .O(new_n1269_));
  NAND     g1253(.a(new_n1269_), .b(new_n1267_), .O(new_n1270_));
  AND      g1254(.a(new_n1270_), .b(i_2_1_51_0), .O(new_n1271_));
  OR       g1255(.a(new_n1271_), .b(new_n1266_), .O(new_n1272_));
  OR       g1256(.a(new_n1272_), .b(new_n1264_), .O(new_n1273_));
  AND      g1257(.a(new_n1273_), .b(i_2_1_70_0), .O(new_n1274_));
  AND      g1258(.a(new_n794_), .b(i_2_1_38_0), .O(new_n1275_));
  OR       g1259(.a(new_n470_), .b(new_n358_), .O(new_n1276_));
  OR       g1260(.a(new_n212_), .b(new_n19_), .O(new_n1277_));
  OR       g1261(.a(new_n1277_), .b(new_n1276_), .O(new_n1278_));
  OR       g1262(.a(new_n1278_), .b(new_n1275_), .O(new_n1279_));
  AND      g1263(.a(new_n1279_), .b(i_2_1_41_0), .O(new_n1280_));
  OR       g1264(.a(new_n1239_), .b(new_n490_), .O(new_n1281_));
  OR       g1265(.a(new_n1281_), .b(new_n1280_), .O(new_n1282_));
  AND      g1266(.a(new_n1282_), .b(new_n18_), .O(new_n1283_));
  NOT      g1267(.a(new_n164_), .O(new_n1284_));
  OR       g1268(.a(new_n1284_), .b(new_n82_), .O(new_n1285_));
  AND      g1269(.a(new_n1285_), .b(new_n387_), .O(new_n1286_));
  OR       g1270(.a(new_n960_), .b(new_n710_), .O(new_n1287_));
  AND      g1271(.a(new_n266_), .b(i_2_1_34_0), .O(new_n1288_));
  AND      g1272(.a(new_n1288_), .b(new_n1287_), .O(new_n1289_));
  OR       g1273(.a(new_n1289_), .b(new_n1286_), .O(new_n1290_));
  OR       g1274(.a(new_n1290_), .b(new_n1283_), .O(new_n1291_));
  OR       g1275(.a(new_n1291_), .b(new_n1274_), .O(new_n1292_));
  AND      g1276(.a(new_n1292_), .b(i_2_1_68_0), .O(new_n1293_));
  AND      g1277(.a(i_2_1_136_0), .b(new_n18_), .O(new_n1294_));
  NAND     g1278(.a(new_n1294_), .b(i_2_1_57_0), .O(new_n1295_));
  NAND     g1279(.a(new_n1295_), .b(new_n624_), .O(new_n1296_));
  AND      g1280(.a(new_n1296_), .b(i_2_1_38_0), .O(new_n1297_));
  AND      g1281(.a(i_2_1_70_0), .b(new_n18_), .O(new_n1298_));
  AND      g1282(.a(new_n1298_), .b(new_n54_), .O(new_n1299_));
  OR       g1283(.a(new_n1299_), .b(new_n74_), .O(new_n1300_));
  AND      g1284(.a(new_n1300_), .b(new_n19_), .O(new_n1301_));
  OR       g1285(.a(new_n1301_), .b(new_n1297_), .O(new_n1302_));
  OR       g1286(.a(new_n1266_), .b(new_n82_), .O(new_n1303_));
  AND      g1287(.a(new_n1303_), .b(i_2_1_34_0), .O(new_n1304_));
  NOT      g1288(.a(new_n155_), .O(new_n1305_));
  AND      g1289(.a(i_2_1_57_0), .b(new_n18_), .O(new_n1306_));
  AND      g1290(.a(new_n1306_), .b(new_n1305_), .O(new_n1307_));
  OR       g1291(.a(new_n1307_), .b(i_2_1_41_0), .O(new_n1308_));
  AND      g1292(.a(new_n1308_), .b(new_n123_), .O(new_n1309_));
  OR       g1293(.a(new_n1309_), .b(new_n1304_), .O(new_n1310_));
  OR       g1294(.a(new_n1310_), .b(new_n1302_), .O(new_n1311_));
  AND      g1295(.a(new_n1311_), .b(i_2_1_13_0), .O(new_n1312_));
  AND      g1296(.a(new_n306_), .b(new_n19_), .O(new_n1313_));
  AND      g1297(.a(i_2_1_135_0), .b(new_n18_), .O(new_n1314_));
  OR       g1298(.a(new_n1314_), .b(new_n73_), .O(new_n1315_));
  AND      g1299(.a(new_n1315_), .b(new_n666_), .O(new_n1316_));
  OR       g1300(.a(new_n1316_), .b(new_n1313_), .O(new_n1317_));
  AND      g1301(.a(new_n1317_), .b(i_2_1_41_0), .O(new_n1318_));
  OR       g1302(.a(new_n1318_), .b(new_n542_), .O(new_n1319_));
  AND      g1303(.a(new_n1319_), .b(i_2_1_34_0), .O(new_n1320_));
  AND      g1304(.a(new_n1314_), .b(new_n447_), .O(new_n1321_));
  OR       g1305(.a(i_2_1_57_0), .b(i_2_1_51_0), .O(new_n1322_));
  NAND     g1306(.a(new_n741_), .b(new_n27_), .O(new_n1323_));
  OR       g1307(.a(new_n1323_), .b(new_n1322_), .O(new_n1324_));
  OR       g1308(.a(new_n915_), .b(new_n531_), .O(new_n1325_));
  NAND     g1309(.a(new_n1325_), .b(new_n1324_), .O(new_n1326_));
  AND      g1310(.a(new_n1326_), .b(new_n102_), .O(new_n1327_));
  OR       g1311(.a(new_n1327_), .b(new_n1321_), .O(new_n1328_));
  OR       g1312(.a(new_n1328_), .b(new_n1320_), .O(new_n1329_));
  OR       g1313(.a(new_n1329_), .b(new_n1312_), .O(new_n1330_));
  OR       g1314(.a(new_n1330_), .b(new_n1293_), .O(new_n1331_));
  OR       g1315(.a(new_n1331_), .b(new_n1259_), .O(new_n1332_));
  AND      g1316(.a(new_n1332_), .b(i_2_1_32_0), .O(new_n1333_));
  NOT      g1317(.a(new_n727_), .O(new_n1334_));
  AND      g1318(.a(new_n617_), .b(i_2_1_68_0), .O(new_n1335_));
  OR       g1319(.a(new_n1335_), .b(new_n1334_), .O(new_n1336_));
  AND      g1320(.a(new_n1336_), .b(i_2_1_34_0), .O(new_n1337_));
  AND      g1321(.a(new_n1071_), .b(i_2_1_38_0), .O(new_n1338_));
  OR       g1322(.a(i_2_1_68_0), .b(new_n18_), .O(new_n1339_));
  NAND     g1323(.a(new_n1339_), .b(new_n52_), .O(new_n1340_));
  AND      g1324(.a(new_n1340_), .b(new_n20_), .O(new_n1341_));
  OR       g1325(.a(new_n1341_), .b(new_n1338_), .O(new_n1342_));
  OR       g1326(.a(new_n1342_), .b(new_n1337_), .O(new_n1343_));
  AND      g1327(.a(new_n1343_), .b(i_2_1_13_0), .O(new_n1344_));
  AND      g1328(.a(new_n532_), .b(i_2_1_136_0), .O(new_n1345_));
  AND      g1329(.a(new_n1345_), .b(new_n1052_), .O(new_n1346_));
  OR       g1330(.a(i_2_1_136_0), .b(i_2_1_68_0), .O(new_n1347_));
  OR       g1331(.a(new_n1347_), .b(new_n625_), .O(new_n1348_));
  AND      g1332(.a(i_2_1_68_0), .b(new_n220_), .O(new_n1349_));
  NAND     g1333(.a(new_n1349_), .b(new_n199_), .O(new_n1350_));
  NAND     g1334(.a(new_n1350_), .b(new_n1348_), .O(new_n1351_));
  AND      g1335(.a(i_2_1_47_0), .b(new_n892_), .O(new_n1352_));
  AND      g1336(.a(new_n1352_), .b(new_n1351_), .O(new_n1353_));
  OR       g1337(.a(new_n1353_), .b(new_n1346_), .O(new_n1354_));
  OR       g1338(.a(new_n1354_), .b(new_n1344_), .O(new_n1355_));
  AND      g1339(.a(new_n1347_), .b(new_n727_), .O(new_n1356_));
  OR       g1340(.a(new_n1356_), .b(new_n287_), .O(new_n1357_));
  AND      g1341(.a(new_n1357_), .b(new_n19_), .O(new_n1358_));
  AND      g1342(.a(new_n532_), .b(new_n194_), .O(new_n1359_));
  AND      g1343(.a(new_n741_), .b(new_n20_), .O(new_n1360_));
  OR       g1344(.a(new_n660_), .b(new_n77_), .O(new_n1361_));
  OR       g1345(.a(new_n1361_), .b(new_n1360_), .O(new_n1362_));
  OR       g1346(.a(new_n1362_), .b(new_n1359_), .O(new_n1363_));
  OR       g1347(.a(new_n1363_), .b(new_n1358_), .O(new_n1364_));
  AND      g1348(.a(new_n1364_), .b(new_n18_), .O(new_n1365_));
  AND      g1349(.a(new_n257_), .b(i_2_1_38_0), .O(new_n1366_));
  OR       g1350(.a(new_n1366_), .b(new_n964_), .O(new_n1367_));
  AND      g1351(.a(new_n1367_), .b(i_2_1_68_0), .O(new_n1368_));
  OR       g1352(.a(new_n287_), .b(new_n19_), .O(new_n1369_));
  AND      g1353(.a(new_n1369_), .b(new_n20_), .O(new_n1370_));
  OR       g1354(.a(new_n1370_), .b(new_n1368_), .O(new_n1371_));
  AND      g1355(.a(new_n1371_), .b(i_2_1_34_0), .O(new_n1372_));
  OR       g1356(.a(new_n1372_), .b(new_n1365_), .O(new_n1373_));
  OR       g1357(.a(new_n1373_), .b(new_n1355_), .O(new_n1374_));
  AND      g1358(.a(new_n1374_), .b(i_2_1_70_0), .O(new_n1375_));
  OR       g1359(.a(new_n1294_), .b(i_2_1_41_0), .O(new_n1376_));
  AND      g1360(.a(new_n1376_), .b(i_2_1_34_0), .O(new_n1377_));
  AND      g1361(.a(new_n617_), .b(i_2_1_38_0), .O(new_n1378_));
  NAND     g1362(.a(i_2_1_57_0), .b(i_2_1_51_0), .O(new_n1379_));
  AND      g1363(.a(new_n1379_), .b(new_n750_), .O(new_n1380_));
  OR       g1364(.a(new_n1380_), .b(new_n1276_), .O(new_n1381_));
  OR       g1365(.a(new_n1381_), .b(new_n1378_), .O(new_n1382_));
  OR       g1366(.a(new_n1382_), .b(new_n1377_), .O(new_n1383_));
  AND      g1367(.a(new_n1383_), .b(new_n19_), .O(new_n1384_));
  OR       g1368(.a(i_2_1_41_0), .b(i_2_1_32_0), .O(new_n1385_));
  NOT      g1369(.a(new_n1385_), .O(new_n1386_));
  AND      g1370(.a(new_n1386_), .b(new_n125_), .O(new_n1387_));
  OR       g1371(.a(new_n387_), .b(i_2_1_38_0), .O(new_n1388_));
  AND      g1372(.a(new_n1388_), .b(new_n989_), .O(new_n1389_));
  OR       g1373(.a(new_n1389_), .b(new_n1387_), .O(new_n1390_));
  AND      g1374(.a(new_n1390_), .b(new_n781_), .O(new_n1391_));
  OR       g1375(.a(new_n470_), .b(new_n125_), .O(new_n1392_));
  AND      g1376(.a(new_n1392_), .b(new_n1294_), .O(new_n1393_));
  AND      g1377(.a(new_n20_), .b(i_2_1_41_0), .O(new_n1394_));
  AND      g1378(.a(new_n1394_), .b(new_n1238_), .O(new_n1395_));
  OR       g1379(.a(new_n1395_), .b(new_n1393_), .O(new_n1396_));
  OR       g1380(.a(new_n1396_), .b(new_n1391_), .O(new_n1397_));
  OR       g1381(.a(new_n1397_), .b(new_n1384_), .O(new_n1398_));
  AND      g1382(.a(new_n1398_), .b(i_2_1_68_0), .O(new_n1399_));
  OR       g1383(.a(new_n1294_), .b(new_n19_), .O(new_n1400_));
  AND      g1384(.a(new_n1400_), .b(i_2_1_38_0), .O(new_n1401_));
  NAND     g1385(.a(new_n727_), .b(new_n533_), .O(new_n1402_));
  AND      g1386(.a(new_n1402_), .b(i_2_1_13_0), .O(new_n1403_));
  OR       g1387(.a(new_n1403_), .b(new_n1401_), .O(new_n1404_));
  AND      g1388(.a(new_n1404_), .b(new_n20_), .O(new_n1405_));
  AND      g1389(.a(new_n837_), .b(i_2_1_38_0), .O(new_n1406_));
  AND      g1390(.a(new_n1406_), .b(new_n19_), .O(new_n1407_));
  OR       g1391(.a(new_n1407_), .b(new_n1405_), .O(new_n1408_));
  AND      g1392(.a(new_n1408_), .b(i_2_1_34_0), .O(new_n1409_));
  OR       g1393(.a(i_2_1_51_0), .b(i_2_1_46_0), .O(new_n1410_));
  NOT      g1394(.a(new_n1410_), .O(new_n1411_));
  AND      g1395(.a(new_n1411_), .b(new_n1345_), .O(new_n1412_));
  OR       g1396(.a(new_n1412_), .b(new_n1409_), .O(new_n1413_));
  OR       g1397(.a(new_n1413_), .b(new_n1399_), .O(new_n1414_));
  OR       g1398(.a(new_n1414_), .b(new_n1375_), .O(new_n1415_));
  AND      g1399(.a(new_n1415_), .b(i_2_1_135_0), .O(new_n1416_));
  OR       g1400(.a(new_n229_), .b(new_n77_), .O(new_n1417_));
  OR       g1401(.a(new_n18_), .b(i_2_1_13_0), .O(new_n1418_));
  AND      g1402(.a(new_n1418_), .b(new_n1417_), .O(new_n1419_));
  NAND     g1403(.a(new_n1018_), .b(new_n174_), .O(new_n1420_));
  AND      g1404(.a(new_n1420_), .b(i_2_1_41_0), .O(new_n1421_));
  AND      g1405(.a(new_n93_), .b(i_2_1_34_0), .O(new_n1422_));
  OR       g1406(.a(new_n1422_), .b(new_n261_), .O(new_n1423_));
  AND      g1407(.a(new_n1423_), .b(i_2_1_68_0), .O(new_n1424_));
  OR       g1408(.a(new_n1424_), .b(new_n1421_), .O(new_n1425_));
  OR       g1409(.a(new_n1425_), .b(new_n1419_), .O(new_n1426_));
  AND      g1410(.a(new_n1426_), .b(i_2_1_38_0), .O(new_n1427_));
  OR       g1411(.a(i_2_1_135_0), .b(new_n52_), .O(new_n1428_));
  NAND     g1412(.a(new_n1428_), .b(new_n25_), .O(new_n1429_));
  AND      g1413(.a(new_n1429_), .b(new_n18_), .O(new_n1430_));
  OR       g1414(.a(new_n237_), .b(new_n20_), .O(new_n1431_));
  AND      g1415(.a(new_n1431_), .b(i_2_1_34_0), .O(new_n1432_));
  OR       g1416(.a(new_n1432_), .b(new_n1430_), .O(new_n1433_));
  AND      g1417(.a(new_n1433_), .b(i_2_1_41_0), .O(new_n1434_));
  AND      g1418(.a(new_n237_), .b(new_n20_), .O(new_n1435_));
  OR       g1419(.a(new_n1435_), .b(new_n1434_), .O(new_n1436_));
  AND      g1420(.a(new_n1436_), .b(i_2_1_70_0), .O(new_n1437_));
  OR       g1421(.a(new_n1017_), .b(new_n77_), .O(new_n1438_));
  AND      g1422(.a(new_n1438_), .b(i_2_1_38_0), .O(new_n1439_));
  AND      g1423(.a(new_n215_), .b(new_n93_), .O(new_n1440_));
  OR       g1424(.a(new_n1440_), .b(new_n18_), .O(new_n1441_));
  AND      g1425(.a(i_2_1_70_0), .b(i_2_1_47_0), .O(new_n1442_));
  OR       g1426(.a(new_n1442_), .b(new_n215_), .O(new_n1443_));
  AND      g1427(.a(new_n1443_), .b(i_2_1_41_0), .O(new_n1444_));
  AND      g1428(.a(new_n1444_), .b(new_n1441_), .O(new_n1445_));
  OR       g1429(.a(new_n1445_), .b(new_n1439_), .O(new_n1446_));
  AND      g1430(.a(new_n1446_), .b(i_2_1_136_0), .O(new_n1447_));
  OR       g1431(.a(new_n1422_), .b(i_2_1_41_0), .O(new_n1448_));
  AND      g1432(.a(new_n1448_), .b(i_2_1_68_0), .O(new_n1449_));
  AND      g1433(.a(new_n1431_), .b(new_n18_), .O(new_n1450_));
  OR       g1434(.a(i_2_1_135_0), .b(i_2_1_51_0), .O(new_n1451_));
  NOT      g1435(.a(new_n1451_), .O(new_n1452_));
  AND      g1436(.a(new_n53_), .b(i_2_1_47_0), .O(new_n1453_));
  OR       g1437(.a(new_n1453_), .b(new_n1452_), .O(new_n1454_));
  AND      g1438(.a(new_n1454_), .b(i_2_1_136_0), .O(new_n1455_));
  OR       g1439(.a(new_n1455_), .b(new_n1450_), .O(new_n1456_));
  OR       g1440(.a(new_n1456_), .b(new_n1449_), .O(new_n1457_));
  AND      g1441(.a(new_n1457_), .b(i_2_1_13_0), .O(new_n1458_));
  OR       g1442(.a(new_n1458_), .b(new_n1447_), .O(new_n1459_));
  OR       g1443(.a(new_n1459_), .b(new_n1437_), .O(new_n1460_));
  OR       g1444(.a(new_n1460_), .b(new_n1427_), .O(new_n1461_));
  AND      g1445(.a(new_n1461_), .b(new_n19_), .O(new_n1462_));
  NOT      g1446(.a(new_n1322_), .O(new_n1463_));
  AND      g1447(.a(new_n1463_), .b(new_n231_), .O(new_n1464_));
  AND      g1448(.a(new_n93_), .b(i_2_1_13_0), .O(new_n1465_));
  AND      g1449(.a(new_n1465_), .b(i_2_1_41_0), .O(new_n1466_));
  OR       g1450(.a(new_n1466_), .b(new_n1464_), .O(new_n1467_));
  AND      g1451(.a(new_n1467_), .b(new_n39_), .O(new_n1468_));
  AND      g1452(.a(new_n18_), .b(i_2_1_13_0), .O(new_n1469_));
  OR       g1453(.a(new_n1469_), .b(new_n77_), .O(new_n1470_));
  OR       g1454(.a(new_n373_), .b(new_n18_), .O(new_n1471_));
  AND      g1455(.a(new_n1471_), .b(new_n1470_), .O(new_n1472_));
  AND      g1456(.a(new_n261_), .b(new_n20_), .O(new_n1473_));
  OR       g1457(.a(new_n1473_), .b(new_n1472_), .O(new_n1474_));
  AND      g1458(.a(new_n1474_), .b(i_2_1_41_0), .O(new_n1475_));
  AND      g1459(.a(new_n1386_), .b(new_n199_), .O(new_n1476_));
  AND      g1460(.a(new_n1476_), .b(new_n573_), .O(new_n1477_));
  OR       g1461(.a(new_n1294_), .b(new_n387_), .O(new_n1478_));
  OR       g1462(.a(new_n1478_), .b(new_n1465_), .O(new_n1479_));
  AND      g1463(.a(new_n1479_), .b(i_2_1_68_0), .O(new_n1480_));
  OR       g1464(.a(new_n1480_), .b(new_n1477_), .O(new_n1481_));
  OR       g1465(.a(new_n1481_), .b(new_n1475_), .O(new_n1482_));
  AND      g1466(.a(new_n1482_), .b(i_2_1_38_0), .O(new_n1483_));
  OR       g1467(.a(new_n1483_), .b(new_n1468_), .O(new_n1484_));
  AND      g1468(.a(new_n1484_), .b(i_2_1_34_0), .O(new_n1485_));
  NAND     g1469(.a(new_n661_), .b(new_n46_), .O(new_n1486_));
  AND      g1470(.a(new_n47_), .b(i_2_1_41_0), .O(new_n1487_));
  AND      g1471(.a(new_n1487_), .b(new_n1486_), .O(new_n1488_));
  OR       g1472(.a(new_n1488_), .b(new_n38_), .O(new_n1489_));
  AND      g1473(.a(new_n1489_), .b(new_n1469_), .O(new_n1490_));
  OR       g1474(.a(new_n1490_), .b(new_n1485_), .O(new_n1491_));
  OR       g1475(.a(new_n1491_), .b(new_n1462_), .O(new_n1492_));
  OR       g1476(.a(new_n1492_), .b(new_n1416_), .O(new_n1493_));
  OR       g1477(.a(new_n1493_), .b(new_n1333_), .O(new_n1494_));
  AND      g1478(.a(new_n1494_), .b(new_n63_), .O(new_n1495_));
  OR       g1479(.a(new_n698_), .b(new_n892_), .O(new_n1496_));
  NAND     g1480(.a(new_n127_), .b(new_n19_), .O(new_n1497_));
  AND      g1481(.a(new_n1497_), .b(new_n533_), .O(new_n1498_));
  NAND     g1482(.a(new_n1498_), .b(new_n1496_), .O(new_n1499_));
  AND      g1483(.a(new_n1499_), .b(i_2_1_68_0), .O(new_n1500_));
  OR       g1484(.a(new_n83_), .b(new_n52_), .O(new_n1501_));
  OR       g1485(.a(new_n21_), .b(i_2_1_38_0), .O(new_n1502_));
  AND      g1486(.a(new_n794_), .b(i_2_1_32_0), .O(new_n1503_));
  AND      g1487(.a(new_n1503_), .b(new_n1502_), .O(new_n1504_));
  AND      g1488(.a(new_n1214_), .b(i_2_1_41_0), .O(new_n1505_));
  NAND     g1489(.a(new_n1505_), .b(new_n1504_), .O(new_n1506_));
  NAND     g1490(.a(new_n1506_), .b(new_n1501_), .O(new_n1507_));
  OR       g1491(.a(new_n1507_), .b(new_n1500_), .O(new_n1508_));
  OR       g1492(.a(new_n1215_), .b(new_n493_), .O(new_n1509_));
  NAND     g1493(.a(new_n155_), .b(i_2_1_38_0), .O(new_n1510_));
  NAND     g1494(.a(new_n1510_), .b(new_n1509_), .O(new_n1511_));
  OR       g1495(.a(new_n175_), .b(i_2_1_34_0), .O(new_n1512_));
  AND      g1496(.a(new_n1512_), .b(new_n892_), .O(new_n1513_));
  OR       g1497(.a(new_n1166_), .b(i_2_1_38_0), .O(new_n1514_));
  AND      g1498(.a(new_n1514_), .b(new_n364_), .O(new_n1515_));
  OR       g1499(.a(new_n1515_), .b(new_n1513_), .O(new_n1516_));
  OR       g1500(.a(new_n1516_), .b(new_n1511_), .O(new_n1517_));
  AND      g1501(.a(new_n1517_), .b(i_2_1_13_0), .O(new_n1518_));
  AND      g1502(.a(new_n1406_), .b(new_n1208_), .O(new_n1519_));
  OR       g1503(.a(new_n1519_), .b(new_n1504_), .O(new_n1520_));
  AND      g1504(.a(new_n1520_), .b(new_n19_), .O(new_n1521_));
  OR       g1505(.a(new_n1521_), .b(new_n1518_), .O(new_n1522_));
  OR       g1506(.a(new_n1522_), .b(new_n1508_), .O(new_n1523_));
  AND      g1507(.a(new_n1523_), .b(new_n18_), .O(new_n1524_));
  AND      g1508(.a(new_n493_), .b(i_2_1_13_0), .O(new_n1525_));
  OR       g1509(.a(new_n1525_), .b(new_n969_), .O(new_n1526_));
  AND      g1510(.a(new_n1526_), .b(new_n279_), .O(new_n1527_));
  AND      g1511(.a(new_n272_), .b(new_n19_), .O(new_n1528_));
  AND      g1512(.a(i_2_1_135_0), .b(i_2_1_49_0), .O(new_n1529_));
  AND      g1513(.a(new_n1529_), .b(new_n52_), .O(new_n1530_));
  OR       g1514(.a(new_n1530_), .b(new_n21_), .O(new_n1531_));
  OR       g1515(.a(new_n1531_), .b(new_n1528_), .O(new_n1532_));
  AND      g1516(.a(new_n1532_), .b(i_2_1_38_0), .O(new_n1533_));
  OR       g1517(.a(new_n709_), .b(new_n549_), .O(new_n1534_));
  OR       g1518(.a(new_n1534_), .b(new_n1101_), .O(new_n1535_));
  AND      g1519(.a(new_n1535_), .b(i_2_1_41_0), .O(new_n1536_));
  NAND     g1520(.a(new_n1428_), .b(new_n459_), .O(new_n1537_));
  AND      g1521(.a(new_n1537_), .b(i_2_1_13_0), .O(new_n1538_));
  OR       g1522(.a(new_n1538_), .b(new_n1165_), .O(new_n1539_));
  OR       g1523(.a(new_n1539_), .b(new_n1536_), .O(new_n1540_));
  OR       g1524(.a(new_n1540_), .b(new_n1533_), .O(new_n1541_));
  AND      g1525(.a(new_n1541_), .b(i_2_1_68_0), .O(new_n1542_));
  OR       g1526(.a(new_n1542_), .b(new_n1527_), .O(new_n1543_));
  OR       g1527(.a(new_n1543_), .b(new_n1524_), .O(new_n1544_));
  AND      g1528(.a(new_n1544_), .b(i_2_1_70_0), .O(new_n1545_));
  OR       g1529(.a(new_n1469_), .b(new_n549_), .O(new_n1546_));
  AND      g1530(.a(new_n1546_), .b(new_n741_), .O(new_n1547_));
  OR       g1531(.a(new_n1547_), .b(new_n380_), .O(new_n1548_));
  AND      g1532(.a(new_n1548_), .b(new_n82_), .O(new_n1549_));
  AND      g1533(.a(i_2_1_41_0), .b(new_n52_), .O(new_n1550_));
  AND      g1534(.a(new_n1550_), .b(new_n380_), .O(new_n1551_));
  OR       g1535(.a(new_n1551_), .b(new_n1549_), .O(new_n1552_));
  OR       g1536(.a(new_n1552_), .b(new_n1545_), .O(new_n1553_));
  OR       g1537(.a(new_n1157_), .b(i_2_1_38_0), .O(new_n1554_));
  AND      g1538(.a(new_n1554_), .b(new_n18_), .O(new_n1555_));
  AND      g1539(.a(new_n127_), .b(i_2_1_38_0), .O(new_n1556_));
  OR       g1540(.a(new_n1556_), .b(new_n1385_), .O(new_n1557_));
  AND      g1541(.a(new_n1557_), .b(new_n1502_), .O(new_n1558_));
  OR       g1542(.a(new_n1558_), .b(new_n1555_), .O(new_n1559_));
  AND      g1543(.a(new_n1559_), .b(i_2_1_13_0), .O(new_n1560_));
  OR       g1544(.a(new_n82_), .b(i_2_1_13_0), .O(new_n1561_));
  OR       g1545(.a(i_2_1_38_0), .b(i_2_1_32_0), .O(new_n1562_));
  AND      g1546(.a(new_n1562_), .b(new_n1561_), .O(new_n1563_));
  AND      g1547(.a(new_n164_), .b(new_n220_), .O(new_n1564_));
  NAND     g1548(.a(new_n1452_), .b(new_n893_), .O(new_n1565_));
  NAND     g1549(.a(new_n1565_), .b(new_n1564_), .O(new_n1566_));
  OR       g1550(.a(new_n1566_), .b(new_n1563_), .O(new_n1567_));
  AND      g1551(.a(new_n1567_), .b(new_n19_), .O(new_n1568_));
  OR       g1552(.a(new_n1265_), .b(i_2_1_136_0), .O(new_n1569_));
  AND      g1553(.a(new_n1569_), .b(new_n1260_), .O(new_n1570_));
  OR       g1554(.a(new_n1570_), .b(new_n712_), .O(new_n1571_));
  AND      g1555(.a(new_n1571_), .b(i_2_1_32_0), .O(new_n1572_));
  AND      g1556(.a(new_n1569_), .b(new_n617_), .O(new_n1573_));
  OR       g1557(.a(new_n82_), .b(new_n175_), .O(new_n1574_));
  AND      g1558(.a(new_n1574_), .b(new_n1573_), .O(new_n1575_));
  OR       g1559(.a(new_n1575_), .b(new_n1572_), .O(new_n1576_));
  OR       g1560(.a(new_n1576_), .b(new_n1568_), .O(new_n1577_));
  OR       g1561(.a(new_n1577_), .b(new_n1560_), .O(new_n1578_));
  AND      g1562(.a(new_n1578_), .b(i_2_1_34_0), .O(new_n1579_));
  AND      g1563(.a(new_n549_), .b(i_2_1_47_0), .O(new_n1580_));
  OR       g1564(.a(new_n1573_), .b(new_n903_), .O(new_n1581_));
  AND      g1565(.a(new_n1581_), .b(i_2_1_13_0), .O(new_n1582_));
  OR       g1566(.a(new_n1582_), .b(new_n1580_), .O(new_n1583_));
  AND      g1567(.a(new_n1583_), .b(i_2_1_38_0), .O(new_n1584_));
  OR       g1568(.a(i_2_1_51_0), .b(new_n102_), .O(new_n1585_));
  NOT      g1569(.a(new_n1585_), .O(new_n1586_));
  NAND     g1570(.a(new_n96_), .b(new_n220_), .O(new_n1587_));
  AND      g1571(.a(new_n1587_), .b(new_n1586_), .O(new_n1588_));
  XOR      g1572(.a(i_2_1_136_0), .b(i_2_1_51_0), .O(new_n1589_));
  AND      g1573(.a(new_n1589_), .b(new_n387_), .O(new_n1590_));
  OR       g1574(.a(new_n1590_), .b(new_n1588_), .O(new_n1591_));
  AND      g1575(.a(new_n1591_), .b(i_2_1_32_0), .O(new_n1592_));
  AND      g1576(.a(new_n524_), .b(i_2_1_136_0), .O(new_n1593_));
  OR       g1577(.a(new_n1593_), .b(new_n1469_), .O(new_n1594_));
  AND      g1578(.a(new_n1594_), .b(new_n19_), .O(new_n1595_));
  OR       g1579(.a(new_n1595_), .b(new_n1592_), .O(new_n1596_));
  AND      g1580(.a(new_n1596_), .b(i_2_1_135_0), .O(new_n1597_));
  OR       g1581(.a(new_n1597_), .b(new_n1584_), .O(new_n1598_));
  OR       g1582(.a(new_n1598_), .b(new_n1579_), .O(new_n1599_));
  AND      g1583(.a(new_n1599_), .b(i_2_1_68_0), .O(new_n1600_));
  AND      g1584(.a(new_n1561_), .b(new_n231_), .O(new_n1601_));
  OR       g1585(.a(new_n1601_), .b(new_n19_), .O(new_n1602_));
  AND      g1586(.a(new_n1602_), .b(new_n18_), .O(new_n1603_));
  AND      g1587(.a(new_n445_), .b(new_n54_), .O(new_n1604_));
  OR       g1588(.a(new_n1604_), .b(new_n1603_), .O(new_n1605_));
  AND      g1589(.a(new_n1605_), .b(i_2_1_136_0), .O(new_n1606_));
  OR       g1590(.a(new_n1261_), .b(new_n960_), .O(new_n1607_));
  AND      g1591(.a(new_n800_), .b(new_n19_), .O(new_n1608_));
  OR       g1592(.a(new_n1608_), .b(new_n709_), .O(new_n1609_));
  AND      g1593(.a(new_n1609_), .b(new_n1607_), .O(new_n1610_));
  OR       g1594(.a(new_n1610_), .b(new_n1606_), .O(new_n1611_));
  AND      g1595(.a(new_n1611_), .b(i_2_1_34_0), .O(new_n1612_));
  OR       g1596(.a(new_n636_), .b(i_2_1_13_0), .O(new_n1613_));
  AND      g1597(.a(new_n1613_), .b(i_2_1_41_0), .O(new_n1614_));
  AND      g1598(.a(new_n1556_), .b(new_n963_), .O(new_n1615_));
  OR       g1599(.a(new_n1615_), .b(new_n660_), .O(new_n1616_));
  OR       g1600(.a(new_n1616_), .b(new_n1614_), .O(new_n1617_));
  AND      g1601(.a(new_n1617_), .b(i_2_1_34_0), .O(new_n1618_));
  OR       g1602(.a(new_n1349_), .b(new_n287_), .O(new_n1619_));
  AND      g1603(.a(new_n1619_), .b(i_2_1_13_0), .O(new_n1620_));
  OR       g1604(.a(new_n1428_), .b(new_n27_), .O(new_n1621_));
  OR       g1605(.a(new_n1621_), .b(new_n963_), .O(new_n1622_));
  NAND     g1606(.a(new_n1622_), .b(new_n574_), .O(new_n1623_));
  AND      g1607(.a(new_n1623_), .b(new_n102_), .O(new_n1624_));
  OR       g1608(.a(new_n1624_), .b(new_n1620_), .O(new_n1625_));
  OR       g1609(.a(new_n1625_), .b(new_n1618_), .O(new_n1626_));
  AND      g1610(.a(new_n1626_), .b(i_2_1_70_0), .O(new_n1627_));
  AND      g1611(.a(new_n1265_), .b(new_n847_), .O(new_n1628_));
  AND      g1612(.a(new_n1628_), .b(new_n1401_), .O(new_n1629_));
  OR       g1613(.a(new_n1629_), .b(new_n1627_), .O(new_n1630_));
  OR       g1614(.a(new_n1630_), .b(new_n1612_), .O(new_n1631_));
  AND      g1615(.a(new_n1631_), .b(i_2_1_32_0), .O(new_n1632_));
  OR       g1616(.a(new_n1632_), .b(new_n1600_), .O(new_n1633_));
  OR       g1617(.a(new_n1633_), .b(new_n1553_), .O(new_n1634_));
  AND      g1618(.a(new_n1634_), .b(new_n20_), .O(new_n1635_));
  OR       g1619(.a(new_n1529_), .b(new_n18_), .O(new_n1636_));
  NOT      g1620(.a(new_n1314_), .O(new_n1637_));
  AND      g1621(.a(new_n1637_), .b(i_2_1_41_0), .O(new_n1638_));
  AND      g1622(.a(new_n1638_), .b(new_n1636_), .O(new_n1639_));
  AND      g1623(.a(new_n18_), .b(i_2_1_34_0), .O(new_n1640_));
  AND      g1624(.a(new_n18_), .b(i_2_1_32_0), .O(new_n1641_));
  OR       g1625(.a(new_n1641_), .b(new_n1640_), .O(new_n1642_));
  OR       g1626(.a(new_n1642_), .b(new_n1639_), .O(new_n1643_));
  AND      g1627(.a(new_n1643_), .b(i_2_1_70_0), .O(new_n1644_));
  OR       g1628(.a(new_n74_), .b(new_n18_), .O(new_n1645_));
  AND      g1629(.a(new_n1645_), .b(i_2_1_38_0), .O(new_n1646_));
  NAND     g1630(.a(new_n1074_), .b(new_n54_), .O(new_n1647_));
  AND      g1631(.a(new_n1647_), .b(new_n535_), .O(new_n1648_));
  OR       g1632(.a(new_n1648_), .b(new_n1646_), .O(new_n1649_));
  OR       g1633(.a(new_n1649_), .b(new_n1644_), .O(new_n1650_));
  AND      g1634(.a(new_n1650_), .b(i_2_1_136_0), .O(new_n1651_));
  OR       g1635(.a(new_n750_), .b(new_n346_), .O(new_n1652_));
  AND      g1636(.a(new_n1652_), .b(new_n1157_), .O(new_n1653_));
  AND      g1637(.a(new_n169_), .b(i_2_1_32_0), .O(new_n1654_));
  OR       g1638(.a(new_n1529_), .b(new_n1306_), .O(new_n1655_));
  OR       g1639(.a(new_n1655_), .b(new_n1654_), .O(new_n1656_));
  AND      g1640(.a(new_n1656_), .b(i_2_1_38_0), .O(new_n1657_));
  AND      g1641(.a(new_n1529_), .b(i_2_1_47_0), .O(new_n1658_));
  OR       g1642(.a(new_n1658_), .b(i_2_1_41_0), .O(new_n1659_));
  AND      g1643(.a(new_n1659_), .b(i_2_1_32_0), .O(new_n1660_));
  OR       g1644(.a(new_n1641_), .b(new_n532_), .O(new_n1661_));
  AND      g1645(.a(new_n1661_), .b(i_2_1_34_0), .O(new_n1662_));
  OR       g1646(.a(new_n1662_), .b(new_n1660_), .O(new_n1663_));
  OR       g1647(.a(new_n1663_), .b(new_n1657_), .O(new_n1664_));
  AND      g1648(.a(new_n1664_), .b(i_2_1_70_0), .O(new_n1665_));
  OR       g1649(.a(new_n1665_), .b(new_n1653_), .O(new_n1666_));
  OR       g1650(.a(new_n1666_), .b(new_n1651_), .O(new_n1667_));
  AND      g1651(.a(new_n1667_), .b(i_2_1_68_0), .O(new_n1668_));
  AND      g1652(.a(new_n1640_), .b(new_n1190_), .O(new_n1669_));
  AND      g1653(.a(new_n794_), .b(new_n712_), .O(new_n1670_));
  AND      g1654(.a(new_n524_), .b(i_2_1_57_0), .O(new_n1671_));
  OR       g1655(.a(new_n1529_), .b(new_n212_), .O(new_n1672_));
  OR       g1656(.a(new_n1672_), .b(new_n1671_), .O(new_n1673_));
  AND      g1657(.a(new_n1673_), .b(new_n18_), .O(new_n1674_));
  OR       g1658(.a(new_n1674_), .b(new_n1670_), .O(new_n1675_));
  AND      g1659(.a(new_n1675_), .b(i_2_1_70_0), .O(new_n1676_));
  OR       g1660(.a(new_n1676_), .b(new_n1100_), .O(new_n1677_));
  AND      g1661(.a(new_n1677_), .b(i_2_1_32_0), .O(new_n1678_));
  OR       g1662(.a(i_2_1_136_0), .b(i_2_1_32_0), .O(new_n1679_));
  NOT      g1663(.a(new_n1679_), .O(new_n1680_));
  AND      g1664(.a(new_n1680_), .b(new_n1314_), .O(new_n1681_));
  OR       g1665(.a(new_n123_), .b(new_n18_), .O(new_n1682_));
  AND      g1666(.a(new_n1682_), .b(new_n212_), .O(new_n1683_));
  OR       g1667(.a(new_n1683_), .b(new_n1681_), .O(new_n1684_));
  AND      g1668(.a(new_n1684_), .b(i_2_1_41_0), .O(new_n1685_));
  OR       g1669(.a(new_n1685_), .b(new_n1678_), .O(new_n1686_));
  AND      g1670(.a(new_n1686_), .b(i_2_1_38_0), .O(new_n1687_));
  OR       g1671(.a(new_n1687_), .b(new_n1669_), .O(new_n1688_));
  OR       g1672(.a(new_n1688_), .b(new_n1668_), .O(new_n1689_));
  AND      g1673(.a(new_n1689_), .b(new_n19_), .O(new_n1690_));
  AND      g1674(.a(new_n209_), .b(new_n18_), .O(new_n1691_));
  OR       g1675(.a(new_n1691_), .b(i_2_1_38_0), .O(new_n1692_));
  AND      g1676(.a(new_n1692_), .b(new_n229_), .O(new_n1693_));
  OR       g1677(.a(new_n1298_), .b(i_2_1_135_0), .O(new_n1694_));
  AND      g1678(.a(new_n1694_), .b(i_2_1_41_0), .O(new_n1695_));
  AND      g1679(.a(i_2_1_136_0), .b(new_n52_), .O(new_n1696_));
  OR       g1680(.a(new_n1696_), .b(new_n660_), .O(new_n1697_));
  AND      g1681(.a(new_n1697_), .b(new_n18_), .O(new_n1698_));
  AND      g1682(.a(new_n103_), .b(i_2_1_51_0), .O(new_n1699_));
  OR       g1683(.a(new_n1699_), .b(new_n21_), .O(new_n1700_));
  OR       g1684(.a(new_n1700_), .b(new_n1698_), .O(new_n1701_));
  OR       g1685(.a(new_n1701_), .b(new_n1695_), .O(new_n1702_));
  OR       g1686(.a(new_n1702_), .b(new_n1693_), .O(new_n1703_));
  AND      g1687(.a(new_n1703_), .b(i_2_1_32_0), .O(new_n1704_));
  AND      g1688(.a(new_n68_), .b(i_2_1_135_0), .O(new_n1705_));
  OR       g1689(.a(new_n1705_), .b(new_n1315_), .O(new_n1706_));
  AND      g1690(.a(new_n1706_), .b(i_2_1_34_0), .O(new_n1707_));
  OR       g1691(.a(new_n1707_), .b(new_n374_), .O(new_n1708_));
  AND      g1692(.a(new_n1708_), .b(i_2_1_68_0), .O(new_n1709_));
  AND      g1693(.a(i_2_1_57_0), .b(i_2_1_38_0), .O(new_n1710_));
  OR       g1694(.a(new_n1710_), .b(i_2_1_68_0), .O(new_n1711_));
  AND      g1695(.a(new_n1711_), .b(i_2_1_41_0), .O(new_n1712_));
  OR       g1696(.a(new_n774_), .b(new_n215_), .O(new_n1713_));
  AND      g1697(.a(new_n1713_), .b(i_2_1_136_0), .O(new_n1714_));
  OR       g1698(.a(new_n1714_), .b(new_n1712_), .O(new_n1715_));
  AND      g1699(.a(new_n1715_), .b(i_2_1_34_0), .O(new_n1716_));
  OR       g1700(.a(new_n1323_), .b(new_n619_), .O(new_n1717_));
  NAND     g1701(.a(new_n287_), .b(i_2_1_57_0), .O(new_n1718_));
  NAND     g1702(.a(new_n1718_), .b(new_n1717_), .O(new_n1719_));
  AND      g1703(.a(new_n1719_), .b(new_n892_), .O(new_n1720_));
  OR       g1704(.a(new_n1720_), .b(new_n1716_), .O(new_n1721_));
  OR       g1705(.a(new_n1721_), .b(new_n1709_), .O(new_n1722_));
  OR       g1706(.a(new_n1722_), .b(new_n1704_), .O(new_n1723_));
  AND      g1707(.a(new_n1723_), .b(new_n19_), .O(new_n1724_));
  AND      g1708(.a(new_n1223_), .b(new_n18_), .O(new_n1725_));
  AND      g1709(.a(new_n994_), .b(i_2_1_136_0), .O(new_n1726_));
  AND      g1710(.a(new_n1347_), .b(new_n362_), .O(new_n1727_));
  OR       g1711(.a(new_n1727_), .b(new_n1726_), .O(new_n1728_));
  OR       g1712(.a(new_n1728_), .b(new_n1725_), .O(new_n1729_));
  AND      g1713(.a(new_n1729_), .b(i_2_1_34_0), .O(new_n1730_));
  AND      g1714(.a(new_n1569_), .b(new_n103_), .O(new_n1731_));
  OR       g1715(.a(new_n1294_), .b(new_n74_), .O(new_n1732_));
  AND      g1716(.a(new_n1732_), .b(i_2_1_70_0), .O(new_n1733_));
  OR       g1717(.a(new_n1733_), .b(new_n1731_), .O(new_n1734_));
  OR       g1718(.a(new_n1734_), .b(new_n1730_), .O(new_n1735_));
  AND      g1719(.a(new_n1735_), .b(i_2_1_38_0), .O(new_n1736_));
  AND      g1720(.a(new_n1265_), .b(new_n37_), .O(new_n1737_));
  AND      g1721(.a(new_n1265_), .b(new_n45_), .O(new_n1738_));
  AND      g1722(.a(new_n1335_), .b(new_n22_), .O(new_n1739_));
  OR       g1723(.a(new_n1739_), .b(new_n1738_), .O(new_n1740_));
  AND      g1724(.a(new_n1740_), .b(i_2_1_34_0), .O(new_n1741_));
  OR       g1725(.a(new_n1741_), .b(new_n1737_), .O(new_n1742_));
  OR       g1726(.a(new_n1742_), .b(new_n1736_), .O(new_n1743_));
  AND      g1727(.a(new_n1743_), .b(i_2_1_32_0), .O(new_n1744_));
  AND      g1728(.a(new_n1586_), .b(new_n37_), .O(new_n1745_));
  AND      g1729(.a(new_n1682_), .b(i_2_1_136_0), .O(new_n1746_));
  OR       g1730(.a(new_n1746_), .b(new_n1298_), .O(new_n1747_));
  AND      g1731(.a(new_n1747_), .b(new_n567_), .O(new_n1748_));
  AND      g1732(.a(new_n362_), .b(new_n37_), .O(new_n1749_));
  OR       g1733(.a(new_n1261_), .b(i_2_1_136_0), .O(new_n1750_));
  OR       g1734(.a(new_n1750_), .b(new_n1749_), .O(new_n1751_));
  AND      g1735(.a(new_n568_), .b(i_2_1_38_0), .O(new_n1752_));
  AND      g1736(.a(new_n1752_), .b(new_n1751_), .O(new_n1753_));
  OR       g1737(.a(new_n1753_), .b(new_n1748_), .O(new_n1754_));
  AND      g1738(.a(new_n1754_), .b(i_2_1_34_0), .O(new_n1755_));
  OR       g1739(.a(new_n1755_), .b(new_n1745_), .O(new_n1756_));
  OR       g1740(.a(new_n1756_), .b(new_n1744_), .O(new_n1757_));
  OR       g1741(.a(new_n1757_), .b(new_n1724_), .O(new_n1758_));
  AND      g1742(.a(new_n1758_), .b(i_2_1_13_0), .O(new_n1759_));
  AND      g1743(.a(new_n1166_), .b(new_n37_), .O(new_n1760_));
  AND      g1744(.a(new_n1760_), .b(new_n1640_), .O(new_n1761_));
  AND      g1745(.a(i_2_1_68_0), .b(new_n18_), .O(new_n1762_));
  AND      g1746(.a(new_n1762_), .b(new_n127_), .O(new_n1763_));
  OR       g1747(.a(new_n1585_), .b(new_n218_), .O(new_n1764_));
  NOT      g1748(.a(new_n39_), .O(new_n1765_));
  AND      g1749(.a(new_n661_), .b(new_n1765_), .O(new_n1766_));
  NAND     g1750(.a(new_n1766_), .b(new_n1764_), .O(new_n1767_));
  AND      g1751(.a(new_n1767_), .b(i_2_1_32_0), .O(new_n1768_));
  OR       g1752(.a(new_n1768_), .b(new_n1763_), .O(new_n1769_));
  AND      g1753(.a(new_n1769_), .b(i_2_1_34_0), .O(new_n1770_));
  OR       g1754(.a(new_n1641_), .b(new_n1284_), .O(new_n1771_));
  AND      g1755(.a(new_n1771_), .b(new_n660_), .O(new_n1772_));
  OR       g1756(.a(new_n1772_), .b(new_n1770_), .O(new_n1773_));
  AND      g1757(.a(new_n1773_), .b(i_2_1_70_0), .O(new_n1774_));
  AND      g1758(.a(new_n1762_), .b(i_2_1_136_0), .O(new_n1775_));
  AND      g1759(.a(new_n1775_), .b(new_n279_), .O(new_n1776_));
  OR       g1760(.a(new_n1776_), .b(new_n1774_), .O(new_n1777_));
  AND      g1761(.a(new_n1777_), .b(i_2_1_41_0), .O(new_n1778_));
  OR       g1762(.a(new_n1778_), .b(new_n1761_), .O(new_n1779_));
  OR       g1763(.a(new_n1779_), .b(new_n1759_), .O(new_n1780_));
  OR       g1764(.a(new_n1780_), .b(new_n1690_), .O(new_n1781_));
  OR       g1765(.a(new_n1781_), .b(new_n1635_), .O(new_n1782_));
  OR       g1766(.a(new_n1782_), .b(new_n1495_), .O(new_n1783_));
  AND      g1767(.a(new_n1783_), .b(new_n32_), .O(new_n1784_));
  AND      g1768(.a(new_n727_), .b(i_2_1_51_0), .O(new_n1785_));
  NAND     g1769(.a(new_n1785_), .b(new_n399_), .O(new_n1786_));
  NAND     g1770(.a(new_n567_), .b(new_n65_), .O(new_n1787_));
  NAND     g1771(.a(new_n1787_), .b(new_n1002_), .O(new_n1788_));
  OR       g1772(.a(new_n1788_), .b(new_n1786_), .O(new_n1789_));
  XOR      g1773(.a(i_2_1_135_0), .b(new_n20_), .O(new_n1790_));
  AND      g1774(.a(new_n1790_), .b(new_n1564_), .O(new_n1791_));
  OR       g1775(.a(new_n567_), .b(i_2_1_51_0), .O(new_n1792_));
  OR       g1776(.a(new_n1792_), .b(new_n1791_), .O(new_n1793_));
  AND      g1777(.a(new_n1793_), .b(new_n1789_), .O(new_n1794_));
  OR       g1778(.a(new_n128_), .b(new_n21_), .O(new_n1795_));
  OR       g1779(.a(new_n1795_), .b(new_n1794_), .O(new_n1796_));
  AND      g1780(.a(new_n1796_), .b(new_n63_), .O(new_n1797_));
  AND      g1781(.a(new_n1298_), .b(i_2_1_136_0), .O(new_n1798_));
  OR       g1782(.a(new_n278_), .b(new_n39_), .O(new_n1799_));
  OR       g1783(.a(new_n1799_), .b(new_n1266_), .O(new_n1800_));
  OR       g1784(.a(new_n1800_), .b(new_n1335_), .O(new_n1801_));
  AND      g1785(.a(new_n1801_), .b(i_2_1_135_0), .O(new_n1802_));
  OR       g1786(.a(new_n1802_), .b(new_n1798_), .O(new_n1803_));
  AND      g1787(.a(new_n1803_), .b(new_n20_), .O(new_n1804_));
  NAND     g1788(.a(new_n1314_), .b(i_2_1_136_0), .O(new_n1805_));
  NAND     g1789(.a(new_n1805_), .b(new_n1024_), .O(new_n1806_));
  AND      g1790(.a(new_n1806_), .b(i_2_1_68_0), .O(new_n1807_));
  OR       g1791(.a(new_n1807_), .b(new_n1804_), .O(new_n1808_));
  OR       g1792(.a(new_n1808_), .b(new_n1797_), .O(new_n1809_));
  AND      g1793(.a(new_n1809_), .b(i_2_1_34_0), .O(new_n1810_));
  OR       g1794(.a(new_n1379_), .b(new_n26_), .O(new_n1811_));
  OR       g1795(.a(new_n762_), .b(i_2_1_51_0), .O(new_n1812_));
  OR       g1796(.a(new_n1812_), .b(new_n152_), .O(new_n1813_));
  AND      g1797(.a(new_n1813_), .b(new_n1811_), .O(new_n1814_));
  OR       g1798(.a(new_n1814_), .b(new_n17_), .O(new_n1815_));
  OR       g1799(.a(new_n54_), .b(i_2_1_49_0), .O(new_n1816_));
  OR       g1800(.a(new_n330_), .b(new_n1816_), .O(new_n1817_));
  NAND     g1801(.a(new_n1817_), .b(new_n1815_), .O(new_n1818_));
  AND      g1802(.a(new_n1818_), .b(new_n53_), .O(new_n1819_));
  AND      g1803(.a(new_n77_), .b(i_2_1_70_0), .O(new_n1820_));
  OR       g1804(.a(new_n1820_), .b(new_n124_), .O(new_n1821_));
  OR       g1805(.a(new_n1821_), .b(new_n654_), .O(new_n1822_));
  AND      g1806(.a(new_n1822_), .b(new_n63_), .O(new_n1823_));
  NAND     g1807(.a(new_n768_), .b(new_n400_), .O(new_n1824_));
  AND      g1808(.a(new_n1824_), .b(new_n18_), .O(new_n1825_));
  AND      g1809(.a(new_n1694_), .b(i_2_1_34_0), .O(new_n1826_));
  AND      g1810(.a(new_n1266_), .b(i_2_1_70_0), .O(new_n1827_));
  OR       g1811(.a(new_n1827_), .b(new_n131_), .O(new_n1828_));
  OR       g1812(.a(new_n1828_), .b(new_n1826_), .O(new_n1829_));
  OR       g1813(.a(new_n1829_), .b(new_n1825_), .O(new_n1830_));
  OR       g1814(.a(new_n1830_), .b(new_n1823_), .O(new_n1831_));
  OR       g1815(.a(new_n1831_), .b(new_n1819_), .O(new_n1832_));
  AND      g1816(.a(new_n1832_), .b(new_n19_), .O(new_n1833_));
  NAND     g1817(.a(new_n1805_), .b(new_n53_), .O(new_n1834_));
  AND      g1818(.a(new_n1834_), .b(i_2_1_41_0), .O(new_n1835_));
  OR       g1819(.a(new_n1835_), .b(new_n1299_), .O(new_n1836_));
  AND      g1820(.a(new_n1836_), .b(new_n77_), .O(new_n1837_));
  AND      g1821(.a(new_n1463_), .b(i_2_1_135_0), .O(new_n1838_));
  OR       g1822(.a(new_n1838_), .b(new_n573_), .O(new_n1839_));
  AND      g1823(.a(new_n1839_), .b(new_n39_), .O(new_n1840_));
  OR       g1824(.a(new_n1137_), .b(new_n278_), .O(new_n1841_));
  AND      g1825(.a(new_n1841_), .b(new_n18_), .O(new_n1842_));
  AND      g1826(.a(new_n1842_), .b(new_n24_), .O(new_n1843_));
  OR       g1827(.a(new_n1843_), .b(new_n78_), .O(new_n1844_));
  AND      g1828(.a(new_n1844_), .b(i_2_1_41_0), .O(new_n1845_));
  OR       g1829(.a(new_n1845_), .b(new_n1840_), .O(new_n1846_));
  AND      g1830(.a(new_n1846_), .b(new_n63_), .O(new_n1847_));
  OR       g1831(.a(new_n1847_), .b(new_n1837_), .O(new_n1848_));
  OR       g1832(.a(new_n1848_), .b(new_n1833_), .O(new_n1849_));
  OR       g1833(.a(new_n1849_), .b(new_n1810_), .O(new_n1850_));
  AND      g1834(.a(new_n1850_), .b(i_2_1_32_0), .O(new_n1851_));
  NAND     g1835(.a(new_n400_), .b(new_n52_), .O(new_n1852_));
  AND      g1836(.a(new_n1852_), .b(new_n65_), .O(new_n1853_));
  OR       g1837(.a(new_n1294_), .b(new_n968_), .O(new_n1854_));
  OR       g1838(.a(new_n1854_), .b(new_n1853_), .O(new_n1855_));
  AND      g1839(.a(new_n1855_), .b(i_2_1_41_0), .O(new_n1856_));
  AND      g1840(.a(new_n1042_), .b(i_2_1_34_0), .O(new_n1857_));
  OR       g1841(.a(new_n1857_), .b(new_n1165_), .O(new_n1858_));
  OR       g1842(.a(new_n1858_), .b(new_n1856_), .O(new_n1859_));
  AND      g1843(.a(new_n1859_), .b(i_2_1_68_0), .O(new_n1860_));
  OR       g1844(.a(new_n550_), .b(i_2_1_51_0), .O(new_n1861_));
  NOT      g1845(.a(new_n1640_), .O(new_n1862_));
  OR       g1846(.a(new_n436_), .b(new_n54_), .O(new_n1863_));
  AND      g1847(.a(new_n1863_), .b(new_n1862_), .O(new_n1864_));
  OR       g1848(.a(new_n1864_), .b(i_2_1_41_0), .O(new_n1865_));
  NAND     g1849(.a(new_n1865_), .b(new_n1861_), .O(new_n1866_));
  OR       g1850(.a(new_n1866_), .b(new_n1860_), .O(new_n1867_));
  AND      g1851(.a(new_n1867_), .b(i_2_1_70_0), .O(new_n1868_));
  AND      g1852(.a(new_n1265_), .b(new_n20_), .O(new_n1869_));
  AND      g1853(.a(new_n257_), .b(new_n74_), .O(new_n1870_));
  OR       g1854(.a(new_n1870_), .b(new_n1869_), .O(new_n1871_));
  AND      g1855(.a(new_n1871_), .b(i_2_1_136_0), .O(new_n1872_));
  OR       g1856(.a(new_n74_), .b(new_n19_), .O(new_n1873_));
  OR       g1857(.a(new_n797_), .b(new_n18_), .O(new_n1874_));
  AND      g1858(.a(new_n1874_), .b(new_n20_), .O(new_n1875_));
  AND      g1859(.a(new_n1875_), .b(new_n1873_), .O(new_n1876_));
  OR       g1860(.a(new_n1876_), .b(new_n1872_), .O(new_n1877_));
  AND      g1861(.a(new_n1877_), .b(i_2_1_68_0), .O(new_n1878_));
  AND      g1862(.a(new_n1852_), .b(new_n1411_), .O(new_n1879_));
  AND      g1863(.a(new_n1360_), .b(new_n1339_), .O(new_n1880_));
  AND      g1864(.a(new_n1411_), .b(i_2_1_68_0), .O(new_n1881_));
  OR       g1865(.a(new_n1881_), .b(new_n1880_), .O(new_n1882_));
  AND      g1866(.a(new_n1882_), .b(new_n127_), .O(new_n1883_));
  OR       g1867(.a(new_n1883_), .b(new_n1879_), .O(new_n1884_));
  OR       g1868(.a(new_n1884_), .b(new_n1878_), .O(new_n1885_));
  OR       g1869(.a(new_n1885_), .b(new_n1868_), .O(new_n1886_));
  AND      g1870(.a(new_n1886_), .b(new_n63_), .O(new_n1887_));
  OR       g1871(.a(new_n1294_), .b(new_n414_), .O(new_n1888_));
  AND      g1872(.a(new_n1888_), .b(i_2_1_34_0), .O(new_n1889_));
  OR       g1873(.a(new_n1052_), .b(new_n417_), .O(new_n1890_));
  AND      g1874(.a(new_n1890_), .b(new_n1054_), .O(new_n1891_));
  OR       g1875(.a(new_n1891_), .b(new_n1889_), .O(new_n1892_));
  AND      g1876(.a(new_n1892_), .b(i_2_1_68_0), .O(new_n1893_));
  AND      g1877(.a(new_n1681_), .b(new_n19_), .O(new_n1894_));
  OR       g1878(.a(new_n1894_), .b(new_n1893_), .O(new_n1895_));
  AND      g1879(.a(new_n1895_), .b(i_2_1_41_0), .O(new_n1896_));
  NAND     g1880(.a(new_n46_), .b(i_2_1_46_0), .O(new_n1897_));
  NAND     g1881(.a(new_n1897_), .b(new_n18_), .O(new_n1898_));
  NAND     g1882(.a(new_n1898_), .b(new_n401_), .O(new_n1899_));
  AND      g1883(.a(new_n1899_), .b(i_2_1_68_0), .O(new_n1900_));
  AND      g1884(.a(new_n124_), .b(new_n18_), .O(new_n1901_));
  OR       g1885(.a(new_n1901_), .b(new_n1900_), .O(new_n1902_));
  AND      g1886(.a(new_n1902_), .b(i_2_1_34_0), .O(new_n1903_));
  AND      g1887(.a(new_n278_), .b(new_n77_), .O(new_n1904_));
  AND      g1888(.a(new_n1904_), .b(new_n1400_), .O(new_n1905_));
  OR       g1889(.a(new_n1905_), .b(new_n1903_), .O(new_n1906_));
  OR       g1890(.a(new_n1906_), .b(new_n1896_), .O(new_n1907_));
  OR       g1891(.a(new_n1907_), .b(new_n1887_), .O(new_n1908_));
  OR       g1892(.a(new_n1908_), .b(new_n1851_), .O(new_n1909_));
  AND      g1893(.a(new_n1909_), .b(i_2_1_38_0), .O(new_n1910_));
  OR       g1894(.a(new_n760_), .b(new_n397_), .O(new_n1911_));
  AND      g1895(.a(new_n1911_), .b(i_2_1_32_0), .O(new_n1912_));
  OR       g1896(.a(new_n1165_), .b(new_n456_), .O(new_n1913_));
  OR       g1897(.a(new_n1913_), .b(new_n1912_), .O(new_n1914_));
  AND      g1898(.a(new_n1914_), .b(new_n63_), .O(new_n1915_));
  OR       g1899(.a(new_n1005_), .b(new_n445_), .O(new_n1916_));
  AND      g1900(.a(new_n1916_), .b(new_n892_), .O(new_n1917_));
  AND      g1901(.a(i_2_1_41_0), .b(i_2_1_32_0), .O(new_n1918_));
  OR       g1902(.a(new_n1918_), .b(new_n148_), .O(new_n1919_));
  OR       g1903(.a(new_n1190_), .b(i_2_1_34_0), .O(new_n1920_));
  AND      g1904(.a(new_n1920_), .b(new_n1919_), .O(new_n1921_));
  OR       g1905(.a(new_n1921_), .b(new_n1917_), .O(new_n1922_));
  OR       g1906(.a(new_n1922_), .b(new_n1915_), .O(new_n1923_));
  AND      g1907(.a(new_n1923_), .b(new_n18_), .O(new_n1924_));
  OR       g1908(.a(new_n1157_), .b(new_n141_), .O(new_n1925_));
  OR       g1909(.a(new_n1925_), .b(new_n97_), .O(new_n1926_));
  AND      g1910(.a(new_n1926_), .b(i_2_1_70_0), .O(new_n1927_));
  NAND     g1911(.a(new_n256_), .b(new_n53_), .O(new_n1928_));
  AND      g1912(.a(new_n1928_), .b(i_2_1_136_0), .O(new_n1929_));
  OR       g1913(.a(new_n1157_), .b(new_n324_), .O(new_n1930_));
  OR       g1914(.a(new_n1930_), .b(new_n1929_), .O(new_n1931_));
  AND      g1915(.a(new_n1931_), .b(i_2_1_41_0), .O(new_n1932_));
  OR       g1916(.a(new_n1932_), .b(new_n1927_), .O(new_n1933_));
  AND      g1917(.a(new_n1933_), .b(new_n19_), .O(new_n1934_));
  NOT      g1918(.a(new_n1529_), .O(new_n1935_));
  AND      g1919(.a(new_n1918_), .b(new_n1935_), .O(new_n1936_));
  AND      g1920(.a(new_n1936_), .b(new_n212_), .O(new_n1937_));
  OR       g1921(.a(new_n1937_), .b(new_n1934_), .O(new_n1938_));
  OR       g1922(.a(new_n1938_), .b(new_n1924_), .O(new_n1939_));
  AND      g1923(.a(new_n1939_), .b(i_2_1_68_0), .O(new_n1940_));
  NOT      g1924(.a(new_n47_), .O(new_n1941_));
  AND      g1925(.a(new_n141_), .b(new_n1941_), .O(new_n1942_));
  OR       g1926(.a(new_n1640_), .b(new_n342_), .O(new_n1943_));
  AND      g1927(.a(new_n1943_), .b(new_n102_), .O(new_n1944_));
  OR       g1928(.a(new_n797_), .b(new_n445_), .O(new_n1945_));
  OR       g1929(.a(new_n1945_), .b(new_n1944_), .O(new_n1946_));
  AND      g1930(.a(new_n1946_), .b(i_2_1_32_0), .O(new_n1947_));
  OR       g1931(.a(new_n1947_), .b(new_n1942_), .O(new_n1948_));
  AND      g1932(.a(new_n1948_), .b(i_2_1_135_0), .O(new_n1949_));
  NAND     g1933(.a(new_n1918_), .b(new_n27_), .O(new_n1950_));
  NAND     g1934(.a(new_n1950_), .b(new_n495_), .O(new_n1951_));
  AND      g1935(.a(new_n1951_), .b(new_n1640_), .O(new_n1952_));
  OR       g1936(.a(new_n271_), .b(new_n18_), .O(new_n1953_));
  AND      g1937(.a(new_n1953_), .b(i_2_1_41_0), .O(new_n1954_));
  AND      g1938(.a(new_n1641_), .b(new_n63_), .O(new_n1955_));
  OR       g1939(.a(new_n1955_), .b(new_n1954_), .O(new_n1956_));
  AND      g1940(.a(new_n1956_), .b(new_n19_), .O(new_n1957_));
  OR       g1941(.a(new_n524_), .b(new_n52_), .O(new_n1958_));
  OR       g1942(.a(i_2_1_51_0), .b(i_2_1_49_0), .O(new_n1959_));
  OR       g1943(.a(new_n1959_), .b(new_n54_), .O(new_n1960_));
  OR       g1944(.a(new_n1960_), .b(new_n327_), .O(new_n1961_));
  NAND     g1945(.a(new_n1961_), .b(new_n1958_), .O(new_n1962_));
  OR       g1946(.a(new_n1962_), .b(new_n1957_), .O(new_n1963_));
  AND      g1947(.a(new_n1963_), .b(i_2_1_136_0), .O(new_n1964_));
  OR       g1948(.a(new_n1964_), .b(new_n1952_), .O(new_n1965_));
  OR       g1949(.a(new_n1965_), .b(new_n1949_), .O(new_n1966_));
  AND      g1950(.a(new_n1966_), .b(i_2_1_70_0), .O(new_n1967_));
  OR       g1951(.a(new_n1967_), .b(new_n1940_), .O(new_n1968_));
  AND      g1952(.a(new_n1968_), .b(new_n20_), .O(new_n1969_));
  AND      g1953(.a(new_n1640_), .b(new_n271_), .O(new_n1970_));
  AND      g1954(.a(new_n1953_), .b(new_n227_), .O(new_n1971_));
  AND      g1955(.a(new_n21_), .b(i_2_1_51_0), .O(new_n1972_));
  OR       g1956(.a(new_n1972_), .b(new_n1971_), .O(new_n1973_));
  AND      g1957(.a(new_n1973_), .b(i_2_1_41_0), .O(new_n1974_));
  NAND     g1958(.a(new_n1637_), .b(new_n1295_), .O(new_n1975_));
  AND      g1959(.a(new_n1975_), .b(new_n1015_), .O(new_n1976_));
  NAND     g1960(.a(new_n1442_), .b(new_n1284_), .O(new_n1977_));
  OR       g1961(.a(new_n1428_), .b(new_n53_), .O(new_n1978_));
  NAND     g1962(.a(new_n1978_), .b(new_n1977_), .O(new_n1979_));
  OR       g1963(.a(new_n1979_), .b(new_n1976_), .O(new_n1980_));
  OR       g1964(.a(new_n1980_), .b(new_n1974_), .O(new_n1981_));
  AND      g1965(.a(new_n1981_), .b(i_2_1_32_0), .O(new_n1982_));
  OR       g1966(.a(new_n1982_), .b(new_n1970_), .O(new_n1983_));
  AND      g1967(.a(new_n1983_), .b(i_2_1_68_0), .O(new_n1984_));
  OR       g1968(.a(new_n1284_), .b(new_n38_), .O(new_n1985_));
  NOT      g1969(.a(new_n1209_), .O(new_n1986_));
  NOT      g1970(.a(new_n1959_), .O(new_n1987_));
  AND      g1971(.a(new_n1987_), .b(new_n1986_), .O(new_n1988_));
  AND      g1972(.a(new_n1988_), .b(new_n1985_), .O(new_n1989_));
  AND      g1973(.a(new_n910_), .b(i_2_1_135_0), .O(new_n1990_));
  OR       g1974(.a(new_n1990_), .b(new_n1017_), .O(new_n1991_));
  AND      g1975(.a(new_n1991_), .b(new_n63_), .O(new_n1992_));
  OR       g1976(.a(new_n1992_), .b(new_n243_), .O(new_n1993_));
  OR       g1977(.a(new_n1993_), .b(new_n1989_), .O(new_n1994_));
  AND      g1978(.a(new_n1994_), .b(i_2_1_41_0), .O(new_n1995_));
  AND      g1979(.a(new_n1640_), .b(new_n278_), .O(new_n1996_));
  OR       g1980(.a(new_n1314_), .b(i_2_1_136_0), .O(new_n1997_));
  NAND     g1981(.a(new_n1997_), .b(i_2_1_34_0), .O(new_n1998_));
  AND      g1982(.a(new_n446_), .b(new_n892_), .O(new_n1999_));
  NAND     g1983(.a(new_n750_), .b(new_n63_), .O(new_n2000_));
  OR       g1984(.a(new_n2000_), .b(new_n1999_), .O(new_n2001_));
  NAND     g1985(.a(new_n2001_), .b(new_n1998_), .O(new_n2002_));
  AND      g1986(.a(new_n2002_), .b(new_n20_), .O(new_n2003_));
  OR       g1987(.a(new_n2003_), .b(new_n1996_), .O(new_n2004_));
  OR       g1988(.a(new_n2004_), .b(new_n1995_), .O(new_n2005_));
  OR       g1989(.a(new_n2005_), .b(new_n1984_), .O(new_n2006_));
  AND      g1990(.a(new_n2006_), .b(new_n19_), .O(new_n2007_));
  NAND     g1991(.a(new_n1775_), .b(new_n342_), .O(new_n2008_));
  NOT      g1992(.a(new_n2008_), .O(new_n2009_));
  AND      g1993(.a(new_n2009_), .b(new_n910_), .O(new_n2010_));
  AND      g1994(.a(new_n921_), .b(new_n231_), .O(new_n2011_));
  AND      g1995(.a(new_n2011_), .b(new_n1746_), .O(new_n2012_));
  OR       g1996(.a(new_n2012_), .b(new_n1990_), .O(new_n2013_));
  AND      g1997(.a(new_n2013_), .b(i_2_1_68_0), .O(new_n2014_));
  AND      g1998(.a(new_n1265_), .b(new_n102_), .O(new_n2015_));
  AND      g1999(.a(new_n2015_), .b(new_n910_), .O(new_n2016_));
  OR       g2000(.a(new_n2016_), .b(new_n2014_), .O(new_n2017_));
  AND      g2001(.a(new_n2017_), .b(new_n63_), .O(new_n2018_));
  OR       g2002(.a(new_n2018_), .b(new_n1760_), .O(new_n2019_));
  AND      g2003(.a(new_n2019_), .b(i_2_1_34_0), .O(new_n2020_));
  OR       g2004(.a(new_n2020_), .b(new_n2010_), .O(new_n2021_));
  OR       g2005(.a(new_n2021_), .b(new_n2007_), .O(new_n2022_));
  OR       g2006(.a(new_n2022_), .b(new_n1969_), .O(new_n2023_));
  OR       g2007(.a(new_n2023_), .b(new_n1910_), .O(new_n2024_));
  AND      g2008(.a(new_n2024_), .b(i_2_1_13_0), .O(new_n2025_));
  OR       g2009(.a(new_n563_), .b(i_2_1_136_0), .O(new_n2026_));
  NAND     g2010(.a(new_n2026_), .b(new_n955_), .O(new_n2027_));
  AND      g2011(.a(new_n2027_), .b(i_2_1_135_0), .O(new_n2028_));
  OR       g2012(.a(new_n148_), .b(new_n19_), .O(new_n2029_));
  AND      g2013(.a(new_n2029_), .b(i_2_1_41_0), .O(new_n2030_));
  AND      g2014(.a(new_n2030_), .b(new_n962_), .O(new_n2031_));
  OR       g2015(.a(new_n617_), .b(new_n55_), .O(new_n2032_));
  NAND     g2016(.a(new_n2032_), .b(new_n1118_), .O(new_n2033_));
  OR       g2017(.a(new_n2033_), .b(new_n2031_), .O(new_n2034_));
  AND      g2018(.a(new_n2034_), .b(new_n20_), .O(new_n2035_));
  OR       g2019(.a(new_n2035_), .b(new_n2028_), .O(new_n2036_));
  AND      g2020(.a(new_n2036_), .b(i_2_1_70_0), .O(new_n2037_));
  NAND     g2021(.a(new_n727_), .b(new_n53_), .O(new_n2038_));
  AND      g2022(.a(new_n169_), .b(new_n531_), .O(new_n2039_));
  AND      g2023(.a(new_n2039_), .b(new_n2038_), .O(new_n2040_));
  OR       g2024(.a(new_n436_), .b(i_2_1_41_0), .O(new_n2041_));
  AND      g2025(.a(new_n300_), .b(new_n674_), .O(new_n2042_));
  NAND     g2026(.a(new_n2042_), .b(new_n2041_), .O(new_n2043_));
  OR       g2027(.a(new_n2043_), .b(new_n2040_), .O(new_n2044_));
  AND      g2028(.a(new_n2044_), .b(i_2_1_135_0), .O(new_n2045_));
  OR       g2029(.a(new_n436_), .b(new_n352_), .O(new_n2046_));
  OR       g2030(.a(new_n954_), .b(new_n469_), .O(new_n2047_));
  NAND     g2031(.a(new_n2047_), .b(new_n436_), .O(new_n2048_));
  OR       g2032(.a(new_n2048_), .b(new_n2030_), .O(new_n2049_));
  NAND     g2033(.a(new_n2049_), .b(i_2_1_70_0), .O(new_n2050_));
  NAND     g2034(.a(new_n2050_), .b(new_n2046_), .O(new_n2051_));
  OR       g2035(.a(new_n2051_), .b(new_n2045_), .O(new_n2052_));
  AND      g2036(.a(new_n2052_), .b(new_n18_), .O(new_n2053_));
  OR       g2037(.a(new_n271_), .b(new_n169_), .O(new_n2054_));
  AND      g2038(.a(new_n2054_), .b(new_n445_), .O(new_n2055_));
  OR       g2039(.a(new_n2055_), .b(new_n2053_), .O(new_n2056_));
  OR       g2040(.a(new_n2056_), .b(new_n2037_), .O(new_n2057_));
  AND      g2041(.a(new_n2057_), .b(i_2_1_38_0), .O(new_n2058_));
  OR       g2042(.a(new_n123_), .b(new_n199_), .O(new_n2059_));
  AND      g2043(.a(new_n2059_), .b(new_n18_), .O(new_n2060_));
  AND      g2044(.a(new_n1726_), .b(new_n1209_), .O(new_n2061_));
  OR       g2045(.a(new_n2061_), .b(new_n2060_), .O(new_n2062_));
  AND      g2046(.a(new_n2062_), .b(new_n63_), .O(new_n2063_));
  AND      g2047(.a(new_n256_), .b(new_n129_), .O(new_n2064_));
  OR       g2048(.a(new_n2064_), .b(new_n2063_), .O(new_n2065_));
  AND      g2049(.a(new_n2065_), .b(new_n445_), .O(new_n2066_));
  OR       g2050(.a(new_n2066_), .b(new_n2058_), .O(new_n2067_));
  AND      g2051(.a(new_n2067_), .b(i_2_1_32_0), .O(new_n2068_));
  OR       g2052(.a(new_n1764_), .b(new_n300_), .O(new_n2069_));
  AND      g2053(.a(new_n2064_), .b(new_n1265_), .O(new_n2070_));
  OR       g2054(.a(new_n278_), .b(i_2_1_38_0), .O(new_n2071_));
  AND      g2055(.a(new_n2071_), .b(new_n1838_), .O(new_n2072_));
  NOT      g2056(.a(new_n446_), .O(new_n2073_));
  AND      g2057(.a(new_n1476_), .b(new_n2073_), .O(new_n2074_));
  NAND     g2058(.a(new_n400_), .b(i_2_1_51_0), .O(new_n2075_));
  AND      g2059(.a(new_n2075_), .b(new_n438_), .O(new_n2076_));
  OR       g2060(.a(new_n2076_), .b(new_n2074_), .O(new_n2077_));
  AND      g2061(.a(new_n2077_), .b(i_2_1_38_0), .O(new_n2078_));
  OR       g2062(.a(new_n2078_), .b(new_n2072_), .O(new_n2079_));
  AND      g2063(.a(new_n2079_), .b(new_n63_), .O(new_n2080_));
  OR       g2064(.a(new_n2080_), .b(new_n2070_), .O(new_n2081_));
  NAND     g2065(.a(new_n2081_), .b(new_n19_), .O(new_n2082_));
  NAND     g2066(.a(new_n2082_), .b(new_n2069_), .O(new_n2083_));
  OR       g2067(.a(new_n2083_), .b(new_n2068_), .O(new_n2084_));
  AND      g2068(.a(new_n2084_), .b(i_2_1_68_0), .O(new_n2085_));
  OR       g2069(.a(new_n1974_), .b(new_n1929_), .O(new_n2086_));
  AND      g2070(.a(new_n2086_), .b(new_n18_), .O(new_n2087_));
  OR       g2071(.a(new_n51_), .b(i_2_1_51_0), .O(new_n2088_));
  NAND     g2072(.a(new_n2088_), .b(new_n193_), .O(new_n2089_));
  AND      g2073(.a(new_n2089_), .b(i_2_1_38_0), .O(new_n2090_));
  OR       g2074(.a(new_n51_), .b(new_n148_), .O(new_n2091_));
  AND      g2075(.a(new_n2091_), .b(new_n20_), .O(new_n2092_));
  OR       g2076(.a(new_n2092_), .b(new_n2090_), .O(new_n2093_));
  OR       g2077(.a(new_n2093_), .b(new_n2087_), .O(new_n2094_));
  AND      g2078(.a(new_n2094_), .b(new_n19_), .O(new_n2095_));
  AND      g2079(.a(new_n1463_), .b(i_2_1_70_0), .O(new_n2096_));
  AND      g2080(.a(new_n18_), .b(i_2_1_49_0), .O(new_n2097_));
  OR       g2081(.a(new_n2097_), .b(new_n954_), .O(new_n2098_));
  OR       g2082(.a(i_2_1_70_0), .b(new_n18_), .O(new_n2099_));
  NAND     g2083(.a(new_n2099_), .b(new_n190_), .O(new_n2100_));
  NAND     g2084(.a(new_n2100_), .b(new_n2098_), .O(new_n2101_));
  AND      g2085(.a(new_n2101_), .b(i_2_1_41_0), .O(new_n2102_));
  AND      g2086(.a(new_n278_), .b(i_2_1_54_0), .O(new_n2103_));
  OR       g2087(.a(new_n2103_), .b(new_n2102_), .O(new_n2104_));
  AND      g2088(.a(new_n2104_), .b(i_2_1_38_0), .O(new_n2105_));
  OR       g2089(.a(new_n2105_), .b(new_n2096_), .O(new_n2106_));
  OR       g2090(.a(new_n2106_), .b(new_n2095_), .O(new_n2107_));
  AND      g2091(.a(new_n2107_), .b(i_2_1_32_0), .O(new_n2108_));
  AND      g2092(.a(new_n169_), .b(new_n124_), .O(new_n2109_));
  AND      g2093(.a(new_n819_), .b(new_n305_), .O(new_n2110_));
  OR       g2094(.a(new_n2110_), .b(new_n2109_), .O(new_n2111_));
  AND      g2095(.a(new_n2111_), .b(i_2_1_38_0), .O(new_n2112_));
  AND      g2096(.a(new_n338_), .b(new_n124_), .O(new_n2113_));
  OR       g2097(.a(new_n549_), .b(new_n73_), .O(new_n2114_));
  AND      g2098(.a(new_n2114_), .b(new_n1452_), .O(new_n2115_));
  OR       g2099(.a(new_n2115_), .b(new_n2113_), .O(new_n2116_));
  OR       g2100(.a(new_n2116_), .b(new_n2112_), .O(new_n2117_));
  AND      g2101(.a(new_n2117_), .b(i_2_1_41_0), .O(new_n2118_));
  AND      g2102(.a(i_2_1_70_0), .b(new_n220_), .O(new_n2119_));
  OR       g2103(.a(new_n2119_), .b(new_n19_), .O(new_n2120_));
  AND      g2104(.a(new_n2120_), .b(new_n271_), .O(new_n2121_));
  OR       g2105(.a(new_n2121_), .b(new_n1298_), .O(new_n2122_));
  AND      g2106(.a(new_n2122_), .b(new_n287_), .O(new_n2123_));
  OR       g2107(.a(new_n2123_), .b(new_n2118_), .O(new_n2124_));
  OR       g2108(.a(new_n2124_), .b(new_n2108_), .O(new_n2125_));
  AND      g2109(.a(new_n2125_), .b(i_2_1_68_0), .O(new_n2126_));
  NOT      g2110(.a(new_n77_), .O(new_n2127_));
  OR       g2111(.a(new_n1585_), .b(new_n20_), .O(new_n2128_));
  OR       g2112(.a(new_n2128_), .b(new_n914_), .O(new_n2129_));
  NAND     g2113(.a(new_n2129_), .b(new_n2127_), .O(new_n2130_));
  AND      g2114(.a(new_n2130_), .b(new_n531_), .O(new_n2131_));
  NAND     g2115(.a(new_n1074_), .b(i_2_1_41_0), .O(new_n2132_));
  OR       g2116(.a(new_n2132_), .b(new_n46_), .O(new_n2133_));
  AND      g2117(.a(new_n1959_), .b(new_n337_), .O(new_n2134_));
  NAND     g2118(.a(new_n2134_), .b(new_n2133_), .O(new_n2135_));
  AND      g2119(.a(new_n2135_), .b(i_2_1_38_0), .O(new_n2136_));
  OR       g2120(.a(new_n1322_), .b(new_n495_), .O(new_n2137_));
  NAND     g2121(.a(new_n2137_), .b(new_n2008_), .O(new_n2138_));
  OR       g2122(.a(new_n2138_), .b(new_n2136_), .O(new_n2139_));
  OR       g2123(.a(new_n2139_), .b(new_n2131_), .O(new_n2140_));
  AND      g2124(.a(new_n2140_), .b(i_2_1_70_0), .O(new_n2141_));
  OR       g2125(.a(new_n1959_), .b(new_n46_), .O(new_n2142_));
  OR       g2126(.a(new_n2097_), .b(i_2_1_136_0), .O(new_n2143_));
  AND      g2127(.a(new_n532_), .b(new_n352_), .O(new_n2144_));
  NAND     g2128(.a(new_n2144_), .b(new_n2143_), .O(new_n2145_));
  NAND     g2129(.a(new_n2145_), .b(new_n2142_), .O(new_n2146_));
  AND      g2130(.a(new_n2146_), .b(i_2_1_68_0), .O(new_n2147_));
  OR       g2131(.a(i_2_1_68_0), .b(i_2_1_47_0), .O(new_n2148_));
  AND      g2132(.a(i_2_1_51_0), .b(new_n63_), .O(new_n2149_));
  AND      g2133(.a(new_n2149_), .b(new_n2148_), .O(new_n2150_));
  OR       g2134(.a(new_n2150_), .b(new_n77_), .O(new_n2151_));
  AND      g2135(.a(new_n2151_), .b(i_2_1_136_0), .O(new_n2152_));
  NAND     g2136(.a(new_n672_), .b(new_n25_), .O(new_n2153_));
  AND      g2137(.a(new_n2153_), .b(new_n1463_), .O(new_n2154_));
  OR       g2138(.a(new_n2154_), .b(new_n567_), .O(new_n2155_));
  OR       g2139(.a(new_n2155_), .b(new_n2152_), .O(new_n2156_));
  AND      g2140(.a(new_n2156_), .b(new_n19_), .O(new_n2157_));
  OR       g2141(.a(new_n2157_), .b(new_n2147_), .O(new_n2158_));
  OR       g2142(.a(new_n2158_), .b(new_n2141_), .O(new_n2159_));
  AND      g2143(.a(new_n2159_), .b(i_2_1_135_0), .O(new_n2160_));
  AND      g2144(.a(new_n532_), .b(new_n63_), .O(new_n2161_));
  OR       g2145(.a(new_n1959_), .b(i_2_1_41_0), .O(new_n2162_));
  NOT      g2146(.a(new_n2162_), .O(new_n2163_));
  OR       g2147(.a(new_n750_), .b(new_n438_), .O(new_n2164_));
  OR       g2148(.a(new_n2164_), .b(new_n2163_), .O(new_n2165_));
  AND      g2149(.a(new_n2165_), .b(new_n20_), .O(new_n2166_));
  OR       g2150(.a(new_n2166_), .b(new_n2161_), .O(new_n2167_));
  OR       g2151(.a(new_n781_), .b(new_n63_), .O(new_n2168_));
  AND      g2152(.a(new_n2168_), .b(new_n19_), .O(new_n2169_));
  AND      g2153(.a(new_n2169_), .b(new_n2167_), .O(new_n2170_));
  OR       g2154(.a(new_n2170_), .b(new_n2160_), .O(new_n2171_));
  AND      g2155(.a(new_n2171_), .b(i_2_1_32_0), .O(new_n2172_));
  OR       g2156(.a(new_n1585_), .b(new_n779_), .O(new_n2173_));
  OR       g2157(.a(new_n1345_), .b(new_n18_), .O(new_n2174_));
  AND      g2158(.a(new_n2174_), .b(new_n324_), .O(new_n2175_));
  AND      g2159(.a(new_n1074_), .b(new_n750_), .O(new_n2176_));
  AND      g2160(.a(new_n2176_), .b(new_n33_), .O(new_n2177_));
  OR       g2161(.a(new_n2119_), .b(new_n1265_), .O(new_n2178_));
  AND      g2162(.a(new_n2178_), .b(new_n287_), .O(new_n2179_));
  OR       g2163(.a(new_n2179_), .b(new_n1298_), .O(new_n2180_));
  OR       g2164(.a(new_n2180_), .b(new_n2177_), .O(new_n2181_));
  AND      g2165(.a(new_n2181_), .b(i_2_1_135_0), .O(new_n2182_));
  OR       g2166(.a(new_n2182_), .b(new_n2175_), .O(new_n2183_));
  AND      g2167(.a(new_n2183_), .b(i_2_1_68_0), .O(new_n2184_));
  AND      g2168(.a(new_n227_), .b(new_n21_), .O(new_n2185_));
  AND      g2169(.a(new_n297_), .b(i_2_1_38_0), .O(new_n2186_));
  AND      g2170(.a(new_n2186_), .b(new_n439_), .O(new_n2187_));
  OR       g2171(.a(new_n2187_), .b(new_n2185_), .O(new_n2188_));
  AND      g2172(.a(new_n2188_), .b(i_2_1_68_0), .O(new_n2189_));
  OR       g2173(.a(new_n412_), .b(new_n82_), .O(new_n2190_));
  AND      g2174(.a(new_n672_), .b(new_n892_), .O(new_n2191_));
  AND      g2175(.a(new_n2191_), .b(new_n2190_), .O(new_n2192_));
  AND      g2176(.a(new_n256_), .b(i_2_1_68_0), .O(new_n2193_));
  AND      g2177(.a(new_n2193_), .b(new_n698_), .O(new_n2194_));
  OR       g2178(.a(new_n2194_), .b(new_n2192_), .O(new_n2195_));
  AND      g2179(.a(new_n2195_), .b(new_n18_), .O(new_n2196_));
  XOR      g2180(.a(i_2_1_136_0), .b(i_2_1_70_0), .O(new_n2197_));
  OR       g2181(.a(new_n2197_), .b(new_n1816_), .O(new_n2198_));
  NAND     g2182(.a(new_n306_), .b(i_2_1_68_0), .O(new_n2199_));
  NAND     g2183(.a(new_n2199_), .b(new_n2198_), .O(new_n2200_));
  AND      g2184(.a(new_n2200_), .b(i_2_1_41_0), .O(new_n2201_));
  OR       g2185(.a(new_n2201_), .b(new_n2196_), .O(new_n2202_));
  OR       g2186(.a(new_n2202_), .b(new_n2189_), .O(new_n2203_));
  AND      g2187(.a(new_n2203_), .b(new_n19_), .O(new_n2204_));
  AND      g2188(.a(new_n2161_), .b(new_n54_), .O(new_n2205_));
  AND      g2189(.a(new_n2205_), .b(new_n1798_), .O(new_n2206_));
  OR       g2190(.a(new_n2206_), .b(new_n2204_), .O(new_n2207_));
  OR       g2191(.a(new_n2207_), .b(new_n2184_), .O(new_n2208_));
  NAND     g2192(.a(new_n2208_), .b(new_n20_), .O(new_n2209_));
  NAND     g2193(.a(new_n2209_), .b(new_n2173_), .O(new_n2210_));
  OR       g2194(.a(new_n2210_), .b(new_n2172_), .O(new_n2211_));
  OR       g2195(.a(new_n2211_), .b(new_n2126_), .O(new_n2212_));
  AND      g2196(.a(new_n2212_), .b(i_2_1_34_0), .O(new_n2213_));
  OR       g2197(.a(new_n1960_), .b(new_n193_), .O(new_n2214_));
  AND      g2198(.a(new_n1451_), .b(new_n399_), .O(new_n2215_));
  OR       g2199(.a(new_n1314_), .b(new_n148_), .O(new_n2216_));
  NAND     g2200(.a(new_n2216_), .b(i_2_1_41_0), .O(new_n2217_));
  OR       g2201(.a(new_n2217_), .b(new_n2215_), .O(new_n2218_));
  NAND     g2202(.a(new_n2218_), .b(new_n2214_), .O(new_n2219_));
  AND      g2203(.a(new_n903_), .b(new_n73_), .O(new_n2220_));
  AND      g2204(.a(new_n2220_), .b(new_n2219_), .O(new_n2221_));
  OR       g2205(.a(new_n2221_), .b(new_n2213_), .O(new_n2222_));
  OR       g2206(.a(new_n2222_), .b(new_n2085_), .O(new_n2223_));
  OR       g2207(.a(new_n2223_), .b(new_n2025_), .O(new_n2224_));
  OR       g2208(.a(new_n2224_), .b(new_n1784_), .O(new_n2225_));
  OR       g2209(.a(new_n2225_), .b(new_n1199_), .O(o_2_1_0_0));
endmodule


