module kernel_2_4 ( 
    i_2_4_12_0, i_2_4_18_0, i_2_4_22_0, i_2_4_24_0, i_2_4_37_0, i_2_4_42_0,
    i_2_4_57_0, i_2_4_70_0, i_2_4_73_0, i_2_4_94_0, i_2_4_109_0,
    i_2_4_117_0, i_2_4_122_0, i_2_4_123_0, i_2_4_133_0,
    o_2_4_0_0  );
  input  i_2_4_12_0, i_2_4_18_0, i_2_4_22_0, i_2_4_24_0, i_2_4_37_0,
    i_2_4_42_0, i_2_4_57_0, i_2_4_70_0, i_2_4_73_0, i_2_4_94_0,
    i_2_4_109_0, i_2_4_117_0, i_2_4_122_0, i_2_4_123_0, i_2_4_133_0;
  output o_2_4_0_0;
  assign o_2_4_0_0 = (~i_2_4_123_0 & ((~i_2_4_133_0 & ((i_2_4_57_0 & ((~i_2_4_117_0 & ((~i_2_4_70_0 & ((~i_2_4_22_0 & ((~i_2_4_12_0 & i_2_4_18_0 & ~i_2_4_42_0 & i_2_4_73_0 & i_2_4_94_0) | (i_2_4_12_0 & i_2_4_24_0 & ~i_2_4_37_0 & i_2_4_42_0 & ~i_2_4_73_0 & ~i_2_4_122_0))) | (~i_2_4_42_0 & ((i_2_4_22_0 & ((~i_2_4_12_0 & ((i_2_4_24_0 & i_2_4_94_0 & i_2_4_109_0) | (i_2_4_18_0 & ~i_2_4_24_0 & i_2_4_73_0 & ~i_2_4_109_0))) | (i_2_4_12_0 & ((i_2_4_94_0 & ((i_2_4_24_0 & (~i_2_4_122_0 | (~i_2_4_37_0 & i_2_4_73_0))) | (~i_2_4_24_0 & i_2_4_73_0 & i_2_4_109_0))) | (~i_2_4_37_0 & ~i_2_4_122_0 & (i_2_4_24_0 | i_2_4_109_0)))) | (~i_2_4_37_0 & ((i_2_4_109_0 & (i_2_4_18_0 | (i_2_4_24_0 & ~i_2_4_122_0))) | (i_2_4_73_0 & ~i_2_4_122_0))))) | (i_2_4_73_0 & ((~i_2_4_37_0 & (((i_2_4_18_0 | (i_2_4_12_0 & ~i_2_4_122_0)) & (i_2_4_24_0 | i_2_4_94_0 | i_2_4_109_0)) | (i_2_4_24_0 & i_2_4_109_0 & ~i_2_4_122_0))) | (i_2_4_18_0 & ~i_2_4_122_0 & (i_2_4_24_0 | i_2_4_109_0)))) | (i_2_4_18_0 & ~i_2_4_122_0 & (~i_2_4_37_0 | (i_2_4_12_0 & i_2_4_24_0 & i_2_4_109_0))))) | (i_2_4_18_0 & ((~i_2_4_122_0 & ((i_2_4_24_0 & ((i_2_4_12_0 & i_2_4_73_0 & (i_2_4_94_0 | i_2_4_109_0)) | i_2_4_22_0 | (i_2_4_94_0 & i_2_4_109_0))) | (i_2_4_22_0 & (~i_2_4_37_0 | i_2_4_94_0)) | (~i_2_4_37_0 & (i_2_4_73_0 | (i_2_4_12_0 & i_2_4_109_0))))) | (i_2_4_109_0 & ((i_2_4_12_0 & ((i_2_4_73_0 & i_2_4_94_0) | (i_2_4_24_0 & ~i_2_4_37_0))) | (i_2_4_24_0 & ~i_2_4_37_0 & i_2_4_94_0))))) | (~i_2_4_37_0 & i_2_4_94_0 & ~i_2_4_122_0 & ((i_2_4_24_0 & i_2_4_109_0) | (i_2_4_22_0 & (i_2_4_12_0 | i_2_4_109_0)))))) | (i_2_4_18_0 & ((~i_2_4_42_0 & ((~i_2_4_12_0 & ((i_2_4_24_0 & i_2_4_70_0 & i_2_4_109_0) | (~i_2_4_73_0 & i_2_4_94_0 & ~i_2_4_122_0))) | (i_2_4_94_0 & ((i_2_4_22_0 & (~i_2_4_37_0 | ~i_2_4_122_0)) | (i_2_4_70_0 & ((i_2_4_24_0 & ~i_2_4_37_0) | (i_2_4_73_0 & i_2_4_109_0))) | (i_2_4_12_0 & i_2_4_73_0 & ~i_2_4_122_0))) | ((~i_2_4_37_0 | ~i_2_4_122_0) & ((i_2_4_22_0 & (i_2_4_24_0 | (i_2_4_12_0 & i_2_4_73_0))) | (i_2_4_12_0 & i_2_4_73_0 & (i_2_4_24_0 | i_2_4_109_0)))) | (i_2_4_109_0 & ((i_2_4_22_0 & (~i_2_4_122_0 | (~i_2_4_37_0 & i_2_4_73_0))) | (~i_2_4_37_0 & ~i_2_4_122_0))) | (~i_2_4_37_0 & ~i_2_4_122_0 & (i_2_4_12_0 | i_2_4_24_0)))) | (i_2_4_109_0 & ((i_2_4_94_0 & ((i_2_4_12_0 & (i_2_4_24_0 | i_2_4_122_0)) | (~i_2_4_122_0 & (i_2_4_22_0 | ~i_2_4_37_0)))) | (i_2_4_24_0 & ((~i_2_4_37_0 & ~i_2_4_122_0) | (i_2_4_22_0 & i_2_4_42_0 & i_2_4_73_0))) | (~i_2_4_37_0 & i_2_4_73_0 & ~i_2_4_122_0))) | (~i_2_4_122_0 & ((i_2_4_22_0 & ((~i_2_4_37_0 & i_2_4_73_0) | (i_2_4_24_0 & i_2_4_94_0))) | (~i_2_4_37_0 & i_2_4_73_0 & (i_2_4_12_0 | i_2_4_24_0 | i_2_4_94_0)))))) | (~i_2_4_37_0 & ~i_2_4_122_0 & ((i_2_4_22_0 & ((~i_2_4_42_0 & ((i_2_4_12_0 & (i_2_4_73_0 | (i_2_4_24_0 & i_2_4_109_0))) | (i_2_4_73_0 & i_2_4_94_0) | ((i_2_4_24_0 | i_2_4_109_0) & (i_2_4_73_0 | i_2_4_94_0)))) | (i_2_4_24_0 & i_2_4_94_0 & i_2_4_109_0) | (i_2_4_12_0 & ((i_2_4_94_0 & i_2_4_109_0) | (i_2_4_24_0 & (i_2_4_94_0 | (i_2_4_73_0 & i_2_4_109_0))))))) | (i_2_4_24_0 & ((~i_2_4_42_0 & i_2_4_73_0 & i_2_4_94_0) | (i_2_4_12_0 & i_2_4_109_0 & (i_2_4_94_0 | (~i_2_4_42_0 & i_2_4_73_0))))) | (i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_42_0 & i_2_4_73_0))) | (i_2_4_12_0 & i_2_4_22_0 & i_2_4_24_0 & i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_42_0 & i_2_4_70_0))) | (i_2_4_18_0 & ((i_2_4_22_0 & ((~i_2_4_42_0 & ((i_2_4_109_0 & ((i_2_4_12_0 & ((i_2_4_73_0 & ~i_2_4_122_0) | (~i_2_4_37_0 & i_2_4_70_0))) | (~i_2_4_37_0 & (i_2_4_94_0 | (~i_2_4_70_0 & i_2_4_73_0))) | (~i_2_4_12_0 & i_2_4_24_0 & i_2_4_70_0) | (~i_2_4_70_0 & i_2_4_73_0 & ~i_2_4_122_0))) | (i_2_4_12_0 & (~i_2_4_37_0 | ~i_2_4_122_0) & (i_2_4_94_0 | (i_2_4_73_0 & (i_2_4_24_0 | ~i_2_4_70_0)))) | (~i_2_4_37_0 & ((i_2_4_24_0 & (i_2_4_94_0 | (~i_2_4_70_0 & i_2_4_73_0))) | ~i_2_4_122_0 | (~i_2_4_70_0 & i_2_4_94_0))))) | (i_2_4_109_0 & ((i_2_4_24_0 & ((i_2_4_12_0 & ~i_2_4_122_0 & (~i_2_4_70_0 | i_2_4_73_0)) | (~i_2_4_12_0 & ~i_2_4_70_0 & i_2_4_94_0))) | (~i_2_4_12_0 & ~i_2_4_37_0 & ~i_2_4_122_0))) | (~i_2_4_37_0 & ~i_2_4_122_0 & ((i_2_4_24_0 & (~i_2_4_70_0 | i_2_4_73_0)) | (i_2_4_73_0 & (i_2_4_12_0 | i_2_4_94_0)))))) | (i_2_4_24_0 & ((i_2_4_109_0 & ((~i_2_4_37_0 & ((i_2_4_94_0 & ((~i_2_4_42_0 & i_2_4_73_0) | (~i_2_4_70_0 & ~i_2_4_122_0))) | (~i_2_4_42_0 & (~i_2_4_122_0 | (i_2_4_12_0 & ~i_2_4_70_0))) | (i_2_4_73_0 & ~i_2_4_122_0) | (i_2_4_12_0 & ((~i_2_4_70_0 & ~i_2_4_122_0) | (i_2_4_42_0 & i_2_4_70_0 & i_2_4_73_0))))) | (~i_2_4_70_0 & i_2_4_73_0 & ~i_2_4_122_0 & i_2_4_12_0 & ~i_2_4_42_0))) | (~i_2_4_122_0 & ((~i_2_4_37_0 & ((~i_2_4_42_0 & (i_2_4_12_0 | ~i_2_4_70_0)) | (i_2_4_73_0 & (~i_2_4_70_0 | i_2_4_94_0)))) | (~i_2_4_42_0 & i_2_4_94_0 & (~i_2_4_70_0 | ~i_2_4_73_0)))))) | (~i_2_4_122_0 & ((i_2_4_94_0 & ((~i_2_4_37_0 & ((i_2_4_12_0 & ~i_2_4_70_0) | ((~i_2_4_42_0 | i_2_4_73_0) & (i_2_4_12_0 | ~i_2_4_70_0 | i_2_4_109_0)))) | (i_2_4_12_0 & ~i_2_4_42_0 & ~i_2_4_70_0 & i_2_4_109_0))) | (~i_2_4_37_0 & ((~i_2_4_42_0 & i_2_4_73_0) | (i_2_4_109_0 & ((~i_2_4_70_0 & i_2_4_73_0) | (~i_2_4_42_0 & (i_2_4_12_0 | ~i_2_4_70_0)))))))))) | (~i_2_4_122_0 & ((~i_2_4_37_0 & ((i_2_4_22_0 & ((i_2_4_24_0 & ((i_2_4_109_0 & ((i_2_4_12_0 & (i_2_4_94_0 | (~i_2_4_42_0 & ~i_2_4_70_0))) | (~i_2_4_42_0 & i_2_4_73_0) | (~i_2_4_70_0 & i_2_4_94_0))) | (~i_2_4_42_0 & i_2_4_73_0 & (~i_2_4_70_0 | i_2_4_94_0)))) | (~i_2_4_70_0 & ((~i_2_4_42_0 & i_2_4_73_0 & i_2_4_94_0) | (i_2_4_12_0 & i_2_4_109_0 & (i_2_4_73_0 | i_2_4_94_0)))))) | (~i_2_4_42_0 & ~i_2_4_70_0 & ((i_2_4_24_0 & i_2_4_94_0 & i_2_4_109_0) | (i_2_4_12_0 & i_2_4_73_0 & ((i_2_4_94_0 & i_2_4_109_0) | (i_2_4_24_0 & (i_2_4_94_0 | i_2_4_109_0)))))))) | (i_2_4_22_0 & ~i_2_4_42_0 & i_2_4_70_0 & i_2_4_73_0 & i_2_4_94_0 & i_2_4_109_0 & i_2_4_117_0))))) | (i_2_4_18_0 & ((~i_2_4_117_0 & ((i_2_4_22_0 & ((i_2_4_94_0 & ((~i_2_4_12_0 & ((~i_2_4_42_0 & ~i_2_4_57_0 & i_2_4_109_0) | (i_2_4_24_0 & i_2_4_73_0 & i_2_4_122_0))) | (i_2_4_12_0 & ((i_2_4_24_0 & (~i_2_4_70_0 | i_2_4_109_0)) | (~i_2_4_42_0 & i_2_4_73_0 & ~i_2_4_122_0))) | (~i_2_4_37_0 & (~i_2_4_122_0 | (~i_2_4_70_0 & i_2_4_73_0))) | (~i_2_4_42_0 & ~i_2_4_70_0 & ~i_2_4_122_0))) | (i_2_4_73_0 & ((i_2_4_12_0 & ((i_2_4_24_0 & ((~i_2_4_37_0 & ~i_2_4_70_0) | (~i_2_4_42_0 & ~i_2_4_122_0))) | (~i_2_4_70_0 & i_2_4_109_0 & (i_2_4_42_0 | ~i_2_4_122_0)))) | (~i_2_4_37_0 & ((~i_2_4_42_0 & ~i_2_4_122_0) | (~i_2_4_57_0 & ~i_2_4_70_0 & i_2_4_109_0))))) | (~i_2_4_122_0 & ((i_2_4_24_0 & ((~i_2_4_37_0 & i_2_4_70_0) | (~i_2_4_42_0 & i_2_4_109_0))) | (~i_2_4_37_0 & (i_2_4_12_0 | i_2_4_109_0 | (~i_2_4_42_0 & ~i_2_4_70_0))))))) | (~i_2_4_42_0 & ((i_2_4_12_0 & ((i_2_4_94_0 & ((i_2_4_24_0 & ((i_2_4_70_0 & i_2_4_109_0) | (~i_2_4_70_0 & i_2_4_73_0 & ~i_2_4_122_0))) | (i_2_4_73_0 & ((~i_2_4_37_0 & i_2_4_70_0 & ~i_2_4_109_0) | (~i_2_4_70_0 & i_2_4_109_0 & ~i_2_4_122_0))))) | (~i_2_4_122_0 & ((~i_2_4_37_0 & (i_2_4_73_0 | (~i_2_4_70_0 & i_2_4_109_0))) | (i_2_4_73_0 & i_2_4_109_0 & i_2_4_24_0 & ~i_2_4_70_0))))) | (~i_2_4_37_0 & ((i_2_4_73_0 & i_2_4_109_0 & i_2_4_24_0 & ~i_2_4_70_0) | (~i_2_4_122_0 & (((i_2_4_24_0 | i_2_4_94_0) & (~i_2_4_70_0 | i_2_4_73_0 | i_2_4_109_0)) | (i_2_4_73_0 & (~i_2_4_70_0 | i_2_4_109_0)))))))) | (~i_2_4_37_0 & ((~i_2_4_122_0 & ((i_2_4_24_0 & (i_2_4_94_0 | (~i_2_4_70_0 & i_2_4_73_0 & i_2_4_109_0))) | (i_2_4_73_0 & i_2_4_94_0 & i_2_4_109_0))) | (i_2_4_12_0 & i_2_4_24_0 & i_2_4_94_0))))) | (~i_2_4_122_0 & ((~i_2_4_42_0 & ((i_2_4_24_0 & ((i_2_4_22_0 & ((i_2_4_12_0 & (~i_2_4_37_0 | (~i_2_4_70_0 & i_2_4_94_0))) | (~i_2_4_37_0 & i_2_4_73_0) | (~i_2_4_12_0 & ((i_2_4_70_0 & i_2_4_94_0) | (~i_2_4_94_0 & ~i_2_4_109_0 & ~i_2_4_70_0 & i_2_4_73_0))))) | (~i_2_4_37_0 & ((i_2_4_12_0 & (i_2_4_73_0 | (~i_2_4_70_0 & i_2_4_109_0))) | (i_2_4_73_0 & (~i_2_4_70_0 | i_2_4_94_0 | i_2_4_109_0)))) | (i_2_4_70_0 & i_2_4_73_0 & i_2_4_94_0 & i_2_4_109_0 & i_2_4_117_0))) | (~i_2_4_37_0 & ((i_2_4_73_0 & (((i_2_4_12_0 | i_2_4_109_0) & (i_2_4_22_0 | i_2_4_94_0)) | (i_2_4_12_0 & i_2_4_109_0) | (~i_2_4_70_0 & (i_2_4_94_0 | i_2_4_109_0)))) | (i_2_4_22_0 & (i_2_4_94_0 | (i_2_4_12_0 & i_2_4_109_0))) | (~i_2_4_70_0 & i_2_4_94_0 & i_2_4_109_0))))) | (~i_2_4_70_0 & ((~i_2_4_37_0 & ((i_2_4_22_0 & (i_2_4_73_0 | (~i_2_4_24_0 & i_2_4_109_0))) | (i_2_4_73_0 & ((i_2_4_24_0 & (i_2_4_12_0 | i_2_4_94_0)) | (i_2_4_12_0 & (i_2_4_94_0 | i_2_4_109_0)))))) | (i_2_4_12_0 & i_2_4_22_0 & i_2_4_24_0 & i_2_4_73_0 & ~i_2_4_94_0 & i_2_4_109_0))) | (i_2_4_22_0 & ~i_2_4_37_0 & ((i_2_4_94_0 & i_2_4_109_0) | (i_2_4_24_0 & (i_2_4_94_0 | (i_2_4_73_0 & i_2_4_109_0))))))) | (i_2_4_22_0 & i_2_4_24_0 & ~i_2_4_37_0 & i_2_4_109_0 & ((i_2_4_12_0 & ~i_2_4_70_0) | (~i_2_4_42_0 & i_2_4_94_0))))) | (~i_2_4_37_0 & ~i_2_4_122_0 & ((i_2_4_73_0 & ((i_2_4_22_0 & ((~i_2_4_117_0 & ((i_2_4_24_0 & ((i_2_4_12_0 & (~i_2_4_70_0 | (~i_2_4_42_0 & i_2_4_109_0))) | (~i_2_4_42_0 & i_2_4_94_0) | (~i_2_4_70_0 & ((~i_2_4_94_0 & i_2_4_109_0) | (i_2_4_94_0 & ~i_2_4_109_0))))) | (i_2_4_12_0 & ~i_2_4_42_0 & ~i_2_4_70_0 & (i_2_4_94_0 | i_2_4_109_0)))) | (~i_2_4_42_0 & i_2_4_94_0 & ((i_2_4_12_0 & i_2_4_109_0) | (~i_2_4_70_0 & (i_2_4_24_0 | i_2_4_109_0)))))) | (i_2_4_24_0 & ~i_2_4_42_0 & i_2_4_94_0 & i_2_4_109_0 & (i_2_4_12_0 | (~i_2_4_70_0 & ~i_2_4_117_0))))) | (i_2_4_12_0 & i_2_4_22_0 & i_2_4_24_0 & ~i_2_4_70_0 & i_2_4_94_0 & ~i_2_4_117_0))))) | (i_2_4_18_0 & ((~i_2_4_37_0 & ((i_2_4_22_0 & ((~i_2_4_42_0 & ((~i_2_4_122_0 & (((i_2_4_24_0 | i_2_4_109_0) & ((~i_2_4_12_0 & ~i_2_4_70_0 & i_2_4_94_0) | (i_2_4_57_0 & i_2_4_73_0 & ~i_2_4_117_0))) | (i_2_4_12_0 & ((i_2_4_24_0 & ((i_2_4_70_0 & i_2_4_94_0) | (i_2_4_57_0 & ~i_2_4_117_0))) | (~i_2_4_70_0 & i_2_4_94_0 & ~i_2_4_117_0) | (i_2_4_57_0 & ((i_2_4_73_0 & i_2_4_94_0 & i_2_4_109_0) | (~i_2_4_70_0 & ~i_2_4_117_0 & (i_2_4_73_0 | i_2_4_109_0)))))) | (i_2_4_94_0 & ((i_2_4_24_0 & i_2_4_109_0 & (i_2_4_57_0 | ~i_2_4_117_0)) | (i_2_4_57_0 & i_2_4_73_0 & (~i_2_4_70_0 | ~i_2_4_117_0)))))) | (i_2_4_12_0 & i_2_4_24_0 & ~i_2_4_57_0 & i_2_4_70_0 & i_2_4_109_0 & ~i_2_4_117_0))) | (~i_2_4_122_0 & ((i_2_4_24_0 & ((i_2_4_73_0 & ((i_2_4_12_0 & ((~i_2_4_70_0 & ~i_2_4_117_0) | (i_2_4_57_0 & i_2_4_109_0))) | (~i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_12_0 & ~i_2_4_70_0))) | (i_2_4_57_0 & ((~i_2_4_70_0 & (i_2_4_94_0 | (i_2_4_109_0 & ~i_2_4_117_0))) | (i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_117_0))))) | (i_2_4_109_0 & ((i_2_4_12_0 & ((i_2_4_94_0 & ~i_2_4_117_0) | (i_2_4_57_0 & ~i_2_4_70_0 & i_2_4_73_0 & i_2_4_117_0))) | (i_2_4_94_0 & ~i_2_4_117_0 & i_2_4_57_0 & ~i_2_4_70_0))))) | (i_2_4_12_0 & i_2_4_24_0 & i_2_4_57_0 & ~i_2_4_70_0 & i_2_4_94_0))) | (~i_2_4_122_0 & ((i_2_4_57_0 & ((i_2_4_73_0 & ((~i_2_4_42_0 & ((~i_2_4_117_0 & (((~i_2_4_70_0 | i_2_4_109_0) & ((i_2_4_24_0 & i_2_4_94_0) | (i_2_4_12_0 & (i_2_4_24_0 | i_2_4_94_0)))) | (~i_2_4_70_0 & i_2_4_109_0 & (i_2_4_12_0 | i_2_4_24_0 | i_2_4_94_0)))) | (i_2_4_94_0 & i_2_4_109_0 & i_2_4_24_0 & ~i_2_4_70_0))) | (i_2_4_94_0 & i_2_4_109_0 & i_2_4_12_0 & i_2_4_24_0))) | (i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_117_0 & i_2_4_12_0 & i_2_4_24_0 & ~i_2_4_70_0))) | (i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_117_0 & i_2_4_12_0 & i_2_4_24_0 & i_2_4_73_0))))) | (i_2_4_22_0 & i_2_4_24_0 & ~i_2_4_42_0 & i_2_4_57_0 & ~i_2_4_70_0 & i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_117_0))) | (i_2_4_12_0 & i_2_4_22_0 & i_2_4_24_0 & ~i_2_4_37_0 & ~i_2_4_42_0 & i_2_4_57_0 & ~i_2_4_70_0 & i_2_4_73_0 & i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_117_0 & ~i_2_4_122_0))) | (i_2_4_18_0 & ~i_2_4_122_0 & ((i_2_4_24_0 & ((i_2_4_12_0 & ((i_2_4_57_0 & ((i_2_4_22_0 & ((~i_2_4_42_0 & ((i_2_4_73_0 & ((~i_2_4_37_0 & ((~i_2_4_70_0 & ~i_2_4_109_0) | (i_2_4_109_0 & ~i_2_4_117_0 & ~i_2_4_133_0))) | (i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_133_0))) | (i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_117_0 & ~i_2_4_133_0))) | (~i_2_4_70_0 & i_2_4_94_0 & i_2_4_117_0))) | (i_2_4_94_0 & ~i_2_4_117_0 & ((~i_2_4_22_0 & ~i_2_4_37_0 & i_2_4_70_0 & ~i_2_4_109_0 & i_2_4_133_0) | (~i_2_4_42_0 & i_2_4_73_0 & i_2_4_109_0 & ~i_2_4_133_0))))) | (i_2_4_73_0 & i_2_4_94_0 & i_2_4_109_0 & i_2_4_22_0 & ~i_2_4_37_0 & ~i_2_4_70_0))) | (~i_2_4_133_0 & ((i_2_4_22_0 & ((~i_2_4_70_0 & i_2_4_109_0 & ((~i_2_4_12_0 & ~i_2_4_117_0 & (i_2_4_94_0 | (~i_2_4_42_0 & i_2_4_73_0))) | (~i_2_4_42_0 & i_2_4_94_0 & i_2_4_117_0))) | (~i_2_4_37_0 & ~i_2_4_42_0 & i_2_4_57_0 & i_2_4_73_0 & i_2_4_94_0 & ~i_2_4_117_0))) | (~i_2_4_12_0 & ~i_2_4_42_0 & ~i_2_4_70_0 & i_2_4_73_0 & i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_117_0))))) | (i_2_4_22_0 & ~i_2_4_42_0 & i_2_4_73_0 & ~i_2_4_133_0 & ((i_2_4_12_0 & ((i_2_4_57_0 & ~i_2_4_117_0 & ((~i_2_4_70_0 & i_2_4_94_0) | (~i_2_4_37_0 & i_2_4_109_0 & (~i_2_4_70_0 | i_2_4_94_0)))) | (~i_2_4_70_0 & i_2_4_94_0 & i_2_4_109_0 & i_2_4_117_0))) | (i_2_4_94_0 & i_2_4_109_0 & ~i_2_4_117_0 & i_2_4_57_0 & ~i_2_4_70_0)))));
endmodule
