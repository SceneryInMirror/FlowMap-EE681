// Benchmark "kernel_2_3" written by ABC on Wed May  4 16:42:44 2022

module kernel_2_3 ( 
    i_2_3_29_0, i_2_3_42_0, i_2_3_43_0, i_2_3_47_0, i_2_3_55_0, i_2_3_68_0,
    i_2_3_72_0, i_2_3_77_0, i_2_3_79_0, i_2_3_86_0, i_2_3_91_0, i_2_3_99_0,
    i_2_3_138_0, i_2_3_142_0, i_2_3_143_0,
    o_2_3_0_0  );
  input  i_2_3_29_0, i_2_3_42_0, i_2_3_43_0, i_2_3_47_0, i_2_3_55_0,
    i_2_3_68_0, i_2_3_72_0, i_2_3_77_0, i_2_3_79_0, i_2_3_86_0, i_2_3_91_0,
    i_2_3_99_0, i_2_3_138_0, i_2_3_142_0, i_2_3_143_0;
  output o_2_3_0_0;
  wire new_n17_, new_n18_, new_n19_, new_n20_, new_n21_, new_n22_, new_n23_,
    new_n24_, new_n25_, new_n26_, new_n27_, new_n28_, new_n29_, new_n30_,
    new_n31_, new_n32_, new_n33_, new_n34_, new_n35_, new_n36_, new_n37_,
    new_n38_, new_n39_, new_n40_, new_n41_, new_n42_, new_n43_, new_n44_,
    new_n45_, new_n46_, new_n47_, new_n48_, new_n49_, new_n50_, new_n51_,
    new_n52_, new_n53_, new_n54_, new_n55_, new_n56_, new_n57_, new_n58_,
    new_n59_, new_n60_, new_n61_, new_n62_, new_n63_, new_n64_, new_n65_,
    new_n66_, new_n67_, new_n68_, new_n69_, new_n70_, new_n71_, new_n72_,
    new_n73_, new_n74_, new_n75_, new_n76_, new_n77_, new_n78_, new_n79_,
    new_n80_, new_n81_, new_n82_, new_n83_, new_n84_, new_n85_, new_n86_,
    new_n87_, new_n88_, new_n89_, new_n90_, new_n91_, new_n92_, new_n93_,
    new_n94_, new_n95_, new_n96_, new_n97_, new_n98_, new_n99_, new_n100_,
    new_n101_, new_n102_, new_n103_, new_n104_, new_n105_, new_n106_,
    new_n107_, new_n108_, new_n109_, new_n110_, new_n111_, new_n112_,
    new_n113_, new_n114_, new_n115_, new_n116_, new_n117_, new_n118_,
    new_n119_, new_n120_, new_n121_, new_n122_, new_n123_, new_n124_,
    new_n125_, new_n126_, new_n127_, new_n128_, new_n129_, new_n130_,
    new_n131_, new_n132_, new_n133_, new_n134_, new_n135_, new_n136_,
    new_n137_, new_n138_, new_n139_, new_n140_, new_n141_, new_n142_,
    new_n143_, new_n144_, new_n145_, new_n146_, new_n147_, new_n148_,
    new_n149_, new_n150_, new_n151_, new_n152_, new_n153_, new_n154_,
    new_n155_, new_n156_, new_n157_, new_n158_, new_n159_, new_n160_,
    new_n161_, new_n162_, new_n163_, new_n164_, new_n165_, new_n166_,
    new_n167_, new_n168_, new_n169_, new_n170_, new_n171_, new_n172_,
    new_n173_, new_n174_, new_n175_, new_n176_, new_n177_, new_n178_,
    new_n179_, new_n180_, new_n181_, new_n182_, new_n183_, new_n184_,
    new_n185_, new_n186_, new_n187_, new_n188_, new_n189_, new_n190_,
    new_n191_, new_n192_, new_n193_, new_n194_, new_n195_, new_n196_,
    new_n197_, new_n198_, new_n199_, new_n200_, new_n201_, new_n202_,
    new_n203_, new_n204_, new_n205_, new_n206_, new_n207_, new_n208_,
    new_n209_, new_n210_, new_n211_, new_n212_, new_n213_, new_n214_,
    new_n215_, new_n216_, new_n217_, new_n218_, new_n219_, new_n220_,
    new_n221_, new_n222_, new_n223_, new_n224_, new_n225_, new_n226_,
    new_n227_, new_n228_, new_n229_, new_n230_, new_n231_, new_n232_,
    new_n233_, new_n234_, new_n235_, new_n236_, new_n237_, new_n238_,
    new_n239_, new_n240_, new_n241_, new_n242_, new_n243_, new_n244_,
    new_n245_, new_n246_, new_n247_, new_n248_, new_n249_, new_n250_,
    new_n251_, new_n252_, new_n253_, new_n254_, new_n255_, new_n256_,
    new_n257_, new_n258_, new_n259_, new_n260_, new_n261_, new_n262_,
    new_n263_, new_n264_, new_n265_, new_n266_, new_n267_, new_n268_,
    new_n269_, new_n270_, new_n271_, new_n272_, new_n273_, new_n274_,
    new_n275_, new_n276_, new_n277_, new_n278_, new_n279_, new_n280_,
    new_n281_, new_n282_, new_n283_, new_n284_, new_n285_, new_n286_,
    new_n287_, new_n288_, new_n289_, new_n290_, new_n291_, new_n292_,
    new_n293_, new_n294_, new_n295_, new_n296_, new_n297_, new_n298_,
    new_n299_, new_n300_, new_n301_, new_n302_, new_n303_, new_n304_,
    new_n305_, new_n306_, new_n307_, new_n308_, new_n309_, new_n310_,
    new_n311_, new_n312_, new_n313_, new_n314_, new_n315_, new_n316_,
    new_n317_, new_n318_, new_n319_, new_n320_, new_n321_, new_n322_,
    new_n323_, new_n324_, new_n325_, new_n326_, new_n327_, new_n328_,
    new_n329_, new_n330_, new_n331_, new_n332_, new_n333_, new_n334_,
    new_n335_, new_n336_, new_n337_, new_n338_, new_n339_, new_n340_,
    new_n341_, new_n342_, new_n343_, new_n344_, new_n345_, new_n346_,
    new_n347_, new_n348_, new_n349_, new_n350_, new_n351_, new_n352_,
    new_n353_, new_n354_, new_n355_, new_n356_, new_n357_, new_n358_,
    new_n359_, new_n360_, new_n361_, new_n362_, new_n363_, new_n364_,
    new_n365_, new_n366_, new_n367_, new_n368_, new_n369_, new_n370_,
    new_n371_, new_n372_, new_n373_, new_n374_, new_n375_, new_n376_,
    new_n377_, new_n378_, new_n379_, new_n380_, new_n381_, new_n382_,
    new_n383_, new_n384_, new_n385_, new_n386_, new_n387_, new_n388_,
    new_n389_, new_n390_, new_n391_, new_n392_, new_n393_, new_n394_,
    new_n395_, new_n396_, new_n397_, new_n398_, new_n399_, new_n400_,
    new_n401_, new_n402_, new_n403_, new_n404_, new_n405_, new_n406_,
    new_n407_, new_n408_, new_n409_, new_n410_, new_n411_, new_n412_,
    new_n413_, new_n414_, new_n415_, new_n416_, new_n417_, new_n418_,
    new_n419_, new_n420_, new_n421_, new_n422_, new_n423_, new_n424_,
    new_n425_, new_n426_, new_n427_, new_n428_, new_n429_, new_n430_,
    new_n431_, new_n432_, new_n433_, new_n434_, new_n435_, new_n436_,
    new_n437_, new_n438_, new_n439_, new_n440_, new_n441_, new_n442_,
    new_n443_, new_n444_, new_n445_, new_n446_, new_n447_, new_n448_,
    new_n449_, new_n450_, new_n451_, new_n452_, new_n453_, new_n454_,
    new_n455_, new_n456_, new_n457_, new_n458_, new_n459_, new_n460_,
    new_n461_, new_n462_, new_n463_, new_n464_, new_n465_, new_n466_,
    new_n467_, new_n468_, new_n469_, new_n470_, new_n471_, new_n472_,
    new_n473_, new_n474_, new_n475_, new_n476_, new_n477_, new_n478_,
    new_n479_, new_n480_, new_n481_, new_n482_, new_n483_, new_n484_,
    new_n485_, new_n486_, new_n487_, new_n488_, new_n489_, new_n490_,
    new_n491_, new_n492_, new_n493_, new_n494_, new_n495_, new_n496_,
    new_n497_, new_n498_, new_n499_, new_n500_, new_n501_, new_n502_,
    new_n503_, new_n504_, new_n505_, new_n506_, new_n507_, new_n508_,
    new_n509_, new_n510_, new_n511_, new_n512_, new_n513_, new_n514_,
    new_n515_, new_n516_, new_n517_, new_n518_, new_n519_, new_n520_,
    new_n521_, new_n522_, new_n523_, new_n524_, new_n525_, new_n526_,
    new_n527_, new_n528_, new_n529_, new_n530_, new_n531_, new_n532_,
    new_n533_, new_n534_, new_n535_, new_n536_, new_n537_, new_n538_,
    new_n539_, new_n540_, new_n541_, new_n542_, new_n543_, new_n544_,
    new_n545_, new_n546_, new_n547_, new_n548_, new_n549_, new_n550_,
    new_n551_, new_n552_, new_n553_, new_n554_, new_n555_, new_n556_,
    new_n557_, new_n558_, new_n559_, new_n560_, new_n561_, new_n562_,
    new_n563_, new_n564_, new_n565_, new_n566_, new_n567_, new_n568_,
    new_n569_, new_n570_, new_n571_, new_n572_, new_n573_, new_n574_,
    new_n575_, new_n576_, new_n577_, new_n578_, new_n579_, new_n580_,
    new_n581_, new_n582_, new_n583_, new_n584_, new_n585_, new_n586_,
    new_n587_, new_n588_, new_n589_, new_n590_, new_n591_, new_n592_,
    new_n593_, new_n594_, new_n595_, new_n596_, new_n597_, new_n598_,
    new_n599_, new_n600_, new_n601_, new_n602_, new_n603_, new_n604_,
    new_n605_, new_n606_, new_n607_, new_n608_, new_n609_, new_n610_,
    new_n611_, new_n612_, new_n613_, new_n614_, new_n615_, new_n616_,
    new_n617_, new_n618_, new_n619_, new_n620_, new_n621_, new_n622_,
    new_n623_, new_n624_, new_n625_, new_n626_, new_n627_, new_n628_,
    new_n629_, new_n630_, new_n631_, new_n632_, new_n633_, new_n634_,
    new_n635_, new_n636_, new_n637_, new_n638_, new_n639_, new_n640_,
    new_n641_, new_n642_, new_n643_, new_n644_, new_n645_, new_n646_,
    new_n647_, new_n648_, new_n649_, new_n650_, new_n651_, new_n652_,
    new_n653_, new_n654_, new_n655_, new_n656_, new_n657_, new_n658_,
    new_n659_, new_n660_, new_n661_, new_n662_, new_n663_, new_n664_,
    new_n665_, new_n666_, new_n667_, new_n668_, new_n669_, new_n670_,
    new_n671_, new_n672_, new_n673_, new_n674_, new_n675_, new_n676_,
    new_n677_, new_n678_, new_n679_, new_n680_, new_n681_, new_n682_,
    new_n683_, new_n684_, new_n685_, new_n686_, new_n687_, new_n688_,
    new_n689_, new_n690_, new_n691_, new_n692_, new_n693_, new_n694_,
    new_n695_, new_n696_, new_n697_, new_n698_, new_n699_, new_n700_,
    new_n701_, new_n702_, new_n703_, new_n704_, new_n705_, new_n706_,
    new_n707_, new_n708_, new_n709_, new_n710_, new_n711_, new_n712_,
    new_n713_, new_n714_, new_n715_, new_n716_, new_n717_, new_n718_,
    new_n719_, new_n720_, new_n721_, new_n722_, new_n723_, new_n724_,
    new_n725_, new_n726_, new_n727_, new_n728_, new_n729_, new_n730_,
    new_n731_, new_n732_, new_n733_, new_n734_, new_n735_, new_n736_,
    new_n737_, new_n738_, new_n739_, new_n740_, new_n741_, new_n742_,
    new_n743_, new_n744_, new_n745_, new_n746_, new_n747_, new_n748_,
    new_n749_, new_n750_, new_n751_, new_n752_, new_n753_, new_n754_,
    new_n755_, new_n756_, new_n757_, new_n758_, new_n759_, new_n760_,
    new_n761_, new_n762_, new_n763_, new_n764_, new_n765_, new_n766_,
    new_n767_, new_n768_, new_n769_, new_n770_, new_n771_, new_n772_,
    new_n773_, new_n774_, new_n775_, new_n776_, new_n777_, new_n778_,
    new_n779_, new_n780_, new_n781_, new_n782_, new_n783_, new_n784_,
    new_n785_, new_n786_, new_n787_, new_n788_, new_n789_, new_n790_,
    new_n791_, new_n792_, new_n793_, new_n794_, new_n795_, new_n796_,
    new_n797_, new_n798_, new_n799_, new_n800_, new_n801_, new_n802_,
    new_n803_, new_n804_, new_n805_, new_n806_, new_n807_, new_n808_,
    new_n809_, new_n810_, new_n811_, new_n812_, new_n813_, new_n814_,
    new_n815_, new_n816_, new_n817_, new_n818_, new_n819_, new_n820_,
    new_n821_, new_n822_, new_n823_, new_n824_, new_n825_, new_n826_,
    new_n827_, new_n828_, new_n829_, new_n830_, new_n831_, new_n832_,
    new_n833_, new_n834_, new_n835_, new_n836_, new_n837_, new_n838_,
    new_n839_, new_n840_, new_n841_, new_n842_, new_n843_, new_n844_,
    new_n845_, new_n846_, new_n847_, new_n848_, new_n849_, new_n850_,
    new_n851_, new_n852_, new_n853_, new_n854_, new_n855_, new_n856_,
    new_n857_, new_n858_, new_n859_, new_n860_, new_n861_, new_n862_,
    new_n863_, new_n864_, new_n865_, new_n866_, new_n867_, new_n868_,
    new_n869_, new_n870_, new_n871_, new_n872_, new_n873_, new_n874_,
    new_n875_, new_n876_, new_n877_, new_n878_, new_n879_, new_n880_,
    new_n881_, new_n882_, new_n883_, new_n884_, new_n885_, new_n886_,
    new_n887_, new_n888_, new_n889_, new_n890_, new_n891_, new_n892_,
    new_n893_, new_n894_, new_n895_, new_n896_, new_n897_, new_n898_,
    new_n899_, new_n900_, new_n901_, new_n902_, new_n903_, new_n904_,
    new_n905_, new_n906_, new_n907_, new_n908_, new_n909_, new_n910_,
    new_n911_, new_n912_, new_n913_, new_n914_, new_n915_, new_n916_,
    new_n917_, new_n918_, new_n919_, new_n920_, new_n921_, new_n922_,
    new_n923_, new_n924_, new_n925_, new_n926_, new_n927_, new_n928_,
    new_n929_, new_n930_, new_n931_, new_n932_, new_n933_, new_n934_,
    new_n935_, new_n936_, new_n937_, new_n938_, new_n939_, new_n940_,
    new_n941_, new_n942_, new_n943_, new_n944_, new_n945_, new_n946_,
    new_n947_, new_n948_, new_n949_, new_n950_, new_n951_, new_n952_,
    new_n953_, new_n954_, new_n955_, new_n956_, new_n957_, new_n958_,
    new_n959_, new_n960_, new_n961_, new_n962_, new_n963_, new_n964_,
    new_n965_, new_n966_, new_n967_, new_n968_, new_n969_, new_n970_,
    new_n971_, new_n972_, new_n973_, new_n974_, new_n975_, new_n976_,
    new_n977_, new_n978_, new_n979_, new_n980_, new_n981_, new_n982_,
    new_n983_, new_n984_, new_n985_, new_n986_, new_n987_, new_n988_,
    new_n989_, new_n990_, new_n991_, new_n992_, new_n993_, new_n994_,
    new_n995_, new_n996_, new_n997_, new_n998_, new_n999_, new_n1000_,
    new_n1001_, new_n1002_, new_n1003_, new_n1004_, new_n1005_, new_n1006_,
    new_n1007_, new_n1008_, new_n1009_, new_n1010_, new_n1011_, new_n1012_,
    new_n1013_, new_n1014_, new_n1015_, new_n1016_, new_n1017_, new_n1018_,
    new_n1019_, new_n1020_, new_n1021_, new_n1022_, new_n1023_, new_n1024_,
    new_n1025_, new_n1026_, new_n1027_, new_n1028_, new_n1029_, new_n1030_,
    new_n1031_, new_n1032_, new_n1033_, new_n1034_, new_n1035_, new_n1036_,
    new_n1037_, new_n1038_, new_n1039_, new_n1040_, new_n1041_, new_n1042_,
    new_n1043_, new_n1044_, new_n1045_, new_n1046_, new_n1047_, new_n1048_,
    new_n1049_, new_n1050_, new_n1051_, new_n1052_, new_n1053_, new_n1054_,
    new_n1055_, new_n1056_, new_n1057_, new_n1058_, new_n1059_, new_n1060_,
    new_n1061_, new_n1062_, new_n1063_, new_n1064_, new_n1065_, new_n1066_,
    new_n1067_, new_n1068_, new_n1069_, new_n1070_, new_n1071_, new_n1072_,
    new_n1073_, new_n1074_, new_n1075_, new_n1076_, new_n1077_, new_n1078_,
    new_n1079_, new_n1080_, new_n1081_, new_n1082_, new_n1083_, new_n1084_,
    new_n1085_, new_n1086_, new_n1087_, new_n1088_, new_n1089_, new_n1090_,
    new_n1091_, new_n1092_, new_n1093_, new_n1094_, new_n1095_, new_n1096_,
    new_n1097_, new_n1098_, new_n1099_, new_n1100_, new_n1101_, new_n1102_,
    new_n1103_, new_n1104_, new_n1105_, new_n1106_, new_n1107_, new_n1108_,
    new_n1109_, new_n1110_, new_n1111_, new_n1112_, new_n1113_, new_n1114_,
    new_n1115_, new_n1116_, new_n1117_, new_n1118_, new_n1119_, new_n1120_,
    new_n1121_, new_n1122_, new_n1123_, new_n1124_, new_n1125_, new_n1126_,
    new_n1127_, new_n1128_, new_n1129_, new_n1130_, new_n1131_, new_n1132_,
    new_n1133_, new_n1134_, new_n1135_, new_n1136_, new_n1137_, new_n1138_,
    new_n1139_, new_n1140_, new_n1141_, new_n1142_, new_n1143_, new_n1144_,
    new_n1145_, new_n1146_, new_n1147_, new_n1148_, new_n1149_, new_n1150_,
    new_n1151_, new_n1152_, new_n1153_, new_n1154_, new_n1155_, new_n1156_,
    new_n1157_, new_n1158_, new_n1159_, new_n1160_, new_n1161_, new_n1162_,
    new_n1163_, new_n1164_, new_n1165_, new_n1166_, new_n1167_, new_n1168_,
    new_n1169_, new_n1170_, new_n1171_, new_n1172_, new_n1173_, new_n1174_,
    new_n1175_, new_n1176_, new_n1177_, new_n1178_, new_n1179_, new_n1180_,
    new_n1181_, new_n1182_, new_n1183_, new_n1184_, new_n1185_, new_n1186_,
    new_n1187_, new_n1188_, new_n1189_, new_n1190_, new_n1191_, new_n1192_,
    new_n1193_, new_n1194_, new_n1195_, new_n1196_, new_n1197_, new_n1198_,
    new_n1199_, new_n1200_, new_n1201_, new_n1202_, new_n1203_, new_n1204_,
    new_n1205_, new_n1206_, new_n1207_, new_n1208_, new_n1209_, new_n1210_,
    new_n1211_, new_n1212_, new_n1213_, new_n1214_, new_n1215_, new_n1216_,
    new_n1217_, new_n1218_, new_n1219_, new_n1220_, new_n1221_, new_n1222_,
    new_n1223_, new_n1224_, new_n1225_, new_n1226_, new_n1227_, new_n1228_,
    new_n1229_, new_n1230_, new_n1231_, new_n1232_, new_n1233_, new_n1234_,
    new_n1235_, new_n1236_, new_n1237_, new_n1238_, new_n1239_, new_n1240_,
    new_n1241_, new_n1242_, new_n1243_, new_n1244_, new_n1245_, new_n1246_,
    new_n1247_, new_n1248_, new_n1249_, new_n1250_, new_n1251_, new_n1252_,
    new_n1253_, new_n1254_, new_n1255_, new_n1256_, new_n1257_, new_n1258_,
    new_n1259_, new_n1260_, new_n1261_, new_n1262_, new_n1263_, new_n1264_,
    new_n1265_, new_n1266_, new_n1267_, new_n1268_, new_n1269_, new_n1270_,
    new_n1271_, new_n1272_, new_n1273_, new_n1274_, new_n1275_, new_n1276_,
    new_n1277_, new_n1278_, new_n1279_, new_n1280_, new_n1281_, new_n1282_,
    new_n1283_, new_n1284_, new_n1285_, new_n1286_, new_n1287_, new_n1288_,
    new_n1289_, new_n1290_, new_n1291_, new_n1292_, new_n1293_, new_n1294_,
    new_n1295_, new_n1296_, new_n1297_, new_n1298_, new_n1299_, new_n1300_,
    new_n1301_, new_n1302_, new_n1303_, new_n1304_, new_n1305_, new_n1306_,
    new_n1307_, new_n1308_, new_n1309_, new_n1310_, new_n1311_, new_n1312_,
    new_n1313_, new_n1314_, new_n1315_, new_n1316_, new_n1317_, new_n1318_,
    new_n1319_, new_n1320_, new_n1321_, new_n1322_, new_n1323_, new_n1324_,
    new_n1325_, new_n1326_, new_n1327_, new_n1328_;
  NOT      g0000(.a(i_2_3_142_0), .O(new_n17_));
  NOT      g0001(.a(i_2_3_143_0), .O(new_n18_));
  NOT      g0002(.a(i_2_3_77_0), .O(new_n19_));
  NOT      g0003(.a(i_2_3_138_0), .O(new_n20_));
  NOT      g0004(.a(i_2_3_79_0), .O(new_n21_));
  OR       g0005(.a(i_2_3_86_0), .b(i_2_3_55_0), .O(new_n22_));
  OR       g0006(.a(i_2_3_47_0), .b(i_2_3_43_0), .O(new_n23_));
  NOT      g0007(.a(i_2_3_91_0), .O(new_n24_));
  NOT      g0008(.a(i_2_3_72_0), .O(new_n25_));
  OR       g0009(.a(new_n25_), .b(i_2_3_42_0), .O(new_n26_));
  AND      g0010(.a(new_n26_), .b(new_n24_), .O(new_n27_));
  NAND     g0011(.a(new_n27_), .b(new_n23_), .O(new_n28_));
  AND      g0012(.a(new_n28_), .b(new_n22_), .O(new_n29_));
  AND      g0013(.a(i_2_3_72_0), .b(i_2_3_55_0), .O(new_n30_));
  NOT      g0014(.a(i_2_3_47_0), .O(new_n31_));
  OR       g0015(.a(i_2_3_86_0), .b(new_n31_), .O(new_n32_));
  AND      g0016(.a(new_n32_), .b(new_n30_), .O(new_n33_));
  OR       g0017(.a(i_2_3_43_0), .b(i_2_3_42_0), .O(new_n34_));
  OR       g0018(.a(new_n34_), .b(i_2_3_47_0), .O(new_n35_));
  NOT      g0019(.a(new_n35_), .O(new_n36_));
  OR       g0020(.a(new_n36_), .b(new_n33_), .O(new_n37_));
  OR       g0021(.a(new_n37_), .b(new_n29_), .O(new_n38_));
  AND      g0022(.a(new_n38_), .b(new_n21_), .O(new_n39_));
  NOT      g0023(.a(i_2_3_99_0), .O(new_n40_));
  AND      g0024(.a(new_n40_), .b(i_2_3_86_0), .O(new_n41_));
  AND      g0025(.a(new_n40_), .b(i_2_3_79_0), .O(new_n42_));
  OR       g0026(.a(new_n42_), .b(i_2_3_72_0), .O(new_n43_));
  OR       g0027(.a(i_2_3_99_0), .b(new_n25_), .O(new_n44_));
  AND      g0028(.a(new_n44_), .b(i_2_3_55_0), .O(new_n45_));
  AND      g0029(.a(new_n45_), .b(new_n43_), .O(new_n46_));
  NAND     g0030(.a(new_n46_), .b(new_n41_), .O(new_n47_));
  OR       g0031(.a(new_n26_), .b(i_2_3_79_0), .O(new_n48_));
  NAND     g0032(.a(new_n48_), .b(new_n47_), .O(new_n49_));
  AND      g0033(.a(new_n49_), .b(i_2_3_43_0), .O(new_n50_));
  AND      g0034(.a(i_2_3_91_0), .b(i_2_3_72_0), .O(new_n51_));
  AND      g0035(.a(new_n51_), .b(new_n31_), .O(new_n52_));
  NOT      g0036(.a(i_2_3_42_0), .O(new_n53_));
  AND      g0037(.a(new_n22_), .b(new_n53_), .O(new_n54_));
  OR       g0038(.a(new_n54_), .b(new_n52_), .O(new_n55_));
  AND      g0039(.a(i_2_3_86_0), .b(i_2_3_55_0), .O(new_n56_));
  OR       g0040(.a(i_2_3_91_0), .b(new_n31_), .O(new_n57_));
  OR       g0041(.a(new_n57_), .b(new_n56_), .O(new_n58_));
  AND      g0042(.a(new_n58_), .b(new_n55_), .O(new_n59_));
  OR       g0043(.a(new_n59_), .b(new_n50_), .O(new_n60_));
  OR       g0044(.a(new_n60_), .b(new_n39_), .O(new_n61_));
  AND      g0045(.a(new_n61_), .b(i_2_3_29_0), .O(new_n62_));
  NAND     g0046(.a(i_2_3_79_0), .b(i_2_3_42_0), .O(new_n63_));
  NAND     g0047(.a(new_n56_), .b(i_2_3_91_0), .O(new_n64_));
  NOT      g0048(.a(new_n64_), .O(new_n65_));
  AND      g0049(.a(i_2_3_86_0), .b(i_2_3_72_0), .O(new_n66_));
  AND      g0050(.a(i_2_3_91_0), .b(i_2_3_55_0), .O(new_n67_));
  OR       g0051(.a(new_n67_), .b(new_n66_), .O(new_n68_));
  OR       g0052(.a(i_2_3_79_0), .b(i_2_3_42_0), .O(new_n69_));
  NOT      g0053(.a(new_n69_), .O(new_n70_));
  OR       g0054(.a(i_2_3_91_0), .b(i_2_3_55_0), .O(new_n71_));
  AND      g0055(.a(new_n71_), .b(new_n70_), .O(new_n72_));
  AND      g0056(.a(new_n72_), .b(new_n68_), .O(new_n73_));
  OR       g0057(.a(new_n73_), .b(new_n65_), .O(new_n74_));
  AND      g0058(.a(new_n74_), .b(new_n63_), .O(new_n75_));
  AND      g0059(.a(i_2_3_91_0), .b(new_n21_), .O(new_n76_));
  NOT      g0060(.a(i_2_3_43_0), .O(new_n77_));
  AND      g0061(.a(i_2_3_91_0), .b(new_n77_), .O(new_n78_));
  OR       g0062(.a(new_n78_), .b(new_n70_), .O(new_n79_));
  AND      g0063(.a(new_n79_), .b(i_2_3_72_0), .O(new_n80_));
  OR       g0064(.a(new_n80_), .b(new_n76_), .O(new_n81_));
  AND      g0065(.a(new_n81_), .b(new_n22_), .O(new_n82_));
  AND      g0066(.a(new_n21_), .b(i_2_3_72_0), .O(new_n83_));
  AND      g0067(.a(new_n83_), .b(new_n56_), .O(new_n84_));
  AND      g0068(.a(new_n71_), .b(i_2_3_86_0), .O(new_n85_));
  OR       g0069(.a(new_n85_), .b(new_n76_), .O(new_n86_));
  AND      g0070(.a(new_n86_), .b(new_n53_), .O(new_n87_));
  OR       g0071(.a(new_n87_), .b(new_n84_), .O(new_n88_));
  OR       g0072(.a(new_n88_), .b(new_n82_), .O(new_n89_));
  AND      g0073(.a(new_n89_), .b(new_n31_), .O(new_n90_));
  OR       g0074(.a(new_n90_), .b(new_n75_), .O(new_n91_));
  OR       g0075(.a(new_n91_), .b(new_n62_), .O(new_n92_));
  AND      g0076(.a(new_n92_), .b(new_n20_), .O(new_n93_));
  OR       g0077(.a(i_2_3_138_0), .b(i_2_3_79_0), .O(new_n94_));
  NAND     g0078(.a(new_n94_), .b(new_n25_), .O(new_n95_));
  OR       g0079(.a(i_2_3_79_0), .b(i_2_3_47_0), .O(new_n96_));
  NAND     g0080(.a(new_n96_), .b(i_2_3_138_0), .O(new_n97_));
  AND      g0081(.a(new_n97_), .b(i_2_3_29_0), .O(new_n98_));
  NOT      g0082(.a(i_2_3_86_0), .O(new_n99_));
  OR       g0083(.a(new_n99_), .b(i_2_3_79_0), .O(new_n100_));
  OR       g0084(.a(i_2_3_138_0), .b(i_2_3_47_0), .O(new_n101_));
  NAND     g0085(.a(new_n101_), .b(new_n100_), .O(new_n102_));
  OR       g0086(.a(new_n102_), .b(new_n98_), .O(new_n103_));
  AND      g0087(.a(new_n103_), .b(new_n95_), .O(new_n104_));
  AND      g0088(.a(i_2_3_86_0), .b(i_2_3_29_0), .O(new_n105_));
  AND      g0089(.a(new_n105_), .b(new_n31_), .O(new_n106_));
  OR       g0090(.a(new_n106_), .b(new_n104_), .O(new_n107_));
  AND      g0091(.a(new_n107_), .b(i_2_3_55_0), .O(new_n108_));
  AND      g0092(.a(i_2_3_86_0), .b(new_n31_), .O(new_n109_));
  AND      g0093(.a(new_n20_), .b(i_2_3_29_0), .O(new_n110_));
  OR       g0094(.a(new_n110_), .b(new_n109_), .O(new_n111_));
  AND      g0095(.a(new_n111_), .b(i_2_3_43_0), .O(new_n112_));
  AND      g0096(.a(i_2_3_86_0), .b(i_2_3_79_0), .O(new_n113_));
  AND      g0097(.a(new_n113_), .b(new_n20_), .O(new_n114_));
  OR       g0098(.a(new_n114_), .b(new_n112_), .O(new_n115_));
  AND      g0099(.a(new_n115_), .b(i_2_3_72_0), .O(new_n116_));
  AND      g0100(.a(new_n105_), .b(new_n76_), .O(new_n117_));
  NAND     g0101(.a(new_n32_), .b(i_2_3_91_0), .O(new_n118_));
  OR       g0102(.a(new_n96_), .b(new_n99_), .O(new_n119_));
  NAND     g0103(.a(new_n119_), .b(new_n118_), .O(new_n120_));
  NAND     g0104(.a(new_n94_), .b(i_2_3_47_0), .O(new_n121_));
  AND      g0105(.a(new_n121_), .b(new_n20_), .O(new_n122_));
  AND      g0106(.a(new_n122_), .b(new_n120_), .O(new_n123_));
  OR       g0107(.a(new_n123_), .b(new_n117_), .O(new_n124_));
  OR       g0108(.a(new_n124_), .b(new_n116_), .O(new_n125_));
  OR       g0109(.a(new_n125_), .b(new_n108_), .O(new_n126_));
  AND      g0110(.a(new_n126_), .b(new_n53_), .O(new_n127_));
  NOT      g0111(.a(new_n26_), .O(new_n128_));
  AND      g0112(.a(new_n67_), .b(new_n128_), .O(new_n129_));
  NAND     g0113(.a(new_n105_), .b(i_2_3_91_0), .O(new_n130_));
  OR       g0114(.a(i_2_3_72_0), .b(i_2_3_47_0), .O(new_n131_));
  NOT      g0115(.a(i_2_3_55_0), .O(new_n132_));
  OR       g0116(.a(i_2_3_138_0), .b(new_n132_), .O(new_n133_));
  OR       g0117(.a(new_n133_), .b(new_n131_), .O(new_n134_));
  NAND     g0118(.a(new_n134_), .b(new_n130_), .O(new_n135_));
  AND      g0119(.a(new_n135_), .b(i_2_3_42_0), .O(new_n136_));
  OR       g0120(.a(new_n136_), .b(new_n129_), .O(new_n137_));
  AND      g0121(.a(new_n137_), .b(i_2_3_79_0), .O(new_n138_));
  AND      g0122(.a(new_n22_), .b(new_n21_), .O(new_n139_));
  OR       g0123(.a(new_n51_), .b(new_n20_), .O(new_n140_));
  OR       g0124(.a(new_n140_), .b(new_n139_), .O(new_n141_));
  AND      g0125(.a(new_n53_), .b(i_2_3_29_0), .O(new_n142_));
  AND      g0126(.a(new_n142_), .b(new_n31_), .O(new_n143_));
  AND      g0127(.a(new_n143_), .b(new_n141_), .O(new_n144_));
  OR       g0128(.a(new_n144_), .b(new_n138_), .O(new_n145_));
  AND      g0129(.a(new_n145_), .b(new_n77_), .O(new_n146_));
  OR       g0130(.a(new_n21_), .b(i_2_3_72_0), .O(new_n147_));
  AND      g0131(.a(new_n147_), .b(i_2_3_86_0), .O(new_n148_));
  OR       g0132(.a(new_n148_), .b(new_n33_), .O(new_n149_));
  AND      g0133(.a(new_n149_), .b(new_n20_), .O(new_n150_));
  AND      g0134(.a(new_n120_), .b(i_2_3_55_0), .O(new_n151_));
  OR       g0135(.a(new_n151_), .b(new_n150_), .O(new_n152_));
  AND      g0136(.a(new_n152_), .b(i_2_3_29_0), .O(new_n153_));
  AND      g0137(.a(new_n20_), .b(i_2_3_91_0), .O(new_n154_));
  NOT      g0138(.a(new_n66_), .O(new_n155_));
  OR       g0139(.a(new_n131_), .b(new_n21_), .O(new_n156_));
  NAND     g0140(.a(new_n156_), .b(new_n155_), .O(new_n157_));
  AND      g0141(.a(new_n157_), .b(new_n154_), .O(new_n158_));
  OR       g0142(.a(new_n158_), .b(new_n153_), .O(new_n159_));
  OR       g0143(.a(new_n159_), .b(new_n146_), .O(new_n160_));
  OR       g0144(.a(new_n160_), .b(new_n127_), .O(new_n161_));
  AND      g0145(.a(new_n161_), .b(i_2_3_99_0), .O(new_n162_));
  AND      g0146(.a(new_n65_), .b(new_n31_), .O(new_n163_));
  AND      g0147(.a(new_n163_), .b(i_2_3_29_0), .O(new_n164_));
  OR       g0148(.a(new_n99_), .b(i_2_3_47_0), .O(new_n165_));
  OR       g0149(.a(new_n132_), .b(i_2_3_43_0), .O(new_n166_));
  OR       g0150(.a(new_n166_), .b(i_2_3_79_0), .O(new_n167_));
  NAND     g0151(.a(new_n167_), .b(new_n165_), .O(new_n168_));
  AND      g0152(.a(new_n168_), .b(i_2_3_72_0), .O(new_n169_));
  OR       g0153(.a(i_2_3_55_0), .b(new_n31_), .O(new_n170_));
  AND      g0154(.a(i_2_3_79_0), .b(i_2_3_43_0), .O(new_n171_));
  NOT      g0155(.a(new_n171_), .O(new_n172_));
  AND      g0156(.a(new_n172_), .b(i_2_3_86_0), .O(new_n173_));
  AND      g0157(.a(new_n173_), .b(new_n170_), .O(new_n174_));
  OR       g0158(.a(new_n174_), .b(new_n169_), .O(new_n175_));
  AND      g0159(.a(new_n175_), .b(i_2_3_29_0), .O(new_n176_));
  OR       g0160(.a(new_n83_), .b(i_2_3_55_0), .O(new_n177_));
  AND      g0161(.a(i_2_3_86_0), .b(new_n77_), .O(new_n178_));
  AND      g0162(.a(new_n178_), .b(new_n31_), .O(new_n179_));
  AND      g0163(.a(new_n179_), .b(new_n177_), .O(new_n180_));
  OR       g0164(.a(new_n180_), .b(new_n176_), .O(new_n181_));
  AND      g0165(.a(new_n181_), .b(i_2_3_91_0), .O(new_n182_));
  AND      g0166(.a(i_2_3_55_0), .b(i_2_3_29_0), .O(new_n183_));
  AND      g0167(.a(new_n183_), .b(new_n31_), .O(new_n184_));
  AND      g0168(.a(new_n184_), .b(new_n148_), .O(new_n185_));
  OR       g0169(.a(new_n185_), .b(new_n182_), .O(new_n186_));
  AND      g0170(.a(new_n186_), .b(new_n53_), .O(new_n187_));
  OR       g0171(.a(new_n187_), .b(new_n164_), .O(new_n188_));
  OR       g0172(.a(new_n188_), .b(new_n162_), .O(new_n189_));
  OR       g0173(.a(new_n189_), .b(new_n93_), .O(new_n190_));
  AND      g0174(.a(new_n190_), .b(i_2_3_68_0), .O(new_n191_));
  OR       g0175(.a(i_2_3_79_0), .b(i_2_3_43_0), .O(new_n192_));
  NOT      g0176(.a(new_n192_), .O(new_n193_));
  AND      g0177(.a(new_n193_), .b(i_2_3_72_0), .O(new_n194_));
  AND      g0178(.a(new_n194_), .b(new_n40_), .O(new_n195_));
  AND      g0179(.a(new_n20_), .b(i_2_3_72_0), .O(new_n196_));
  OR       g0180(.a(new_n196_), .b(new_n46_), .O(new_n197_));
  OR       g0181(.a(new_n197_), .b(new_n195_), .O(new_n198_));
  AND      g0182(.a(new_n198_), .b(new_n31_), .O(new_n199_));
  AND      g0183(.a(new_n21_), .b(i_2_3_55_0), .O(new_n200_));
  NAND     g0184(.a(new_n200_), .b(i_2_3_86_0), .O(new_n201_));
  OR       g0185(.a(new_n66_), .b(new_n20_), .O(new_n202_));
  NAND     g0186(.a(new_n202_), .b(new_n31_), .O(new_n203_));
  NAND     g0187(.a(new_n203_), .b(new_n201_), .O(new_n204_));
  AND      g0188(.a(new_n204_), .b(i_2_3_99_0), .O(new_n205_));
  OR       g0189(.a(i_2_3_99_0), .b(new_n21_), .O(new_n206_));
  AND      g0190(.a(new_n206_), .b(new_n20_), .O(new_n207_));
  AND      g0191(.a(new_n207_), .b(new_n22_), .O(new_n208_));
  OR       g0192(.a(new_n208_), .b(new_n205_), .O(new_n209_));
  OR       g0193(.a(new_n209_), .b(new_n199_), .O(new_n210_));
  AND      g0194(.a(new_n210_), .b(i_2_3_91_0), .O(new_n211_));
  AND      g0195(.a(i_2_3_99_0), .b(new_n21_), .O(new_n212_));
  AND      g0196(.a(i_2_3_55_0), .b(new_n31_), .O(new_n213_));
  AND      g0197(.a(new_n213_), .b(i_2_3_86_0), .O(new_n214_));
  AND      g0198(.a(new_n214_), .b(new_n212_), .O(new_n215_));
  OR       g0199(.a(new_n215_), .b(new_n211_), .O(new_n216_));
  AND      g0200(.a(new_n216_), .b(new_n53_), .O(new_n217_));
  AND      g0201(.a(new_n56_), .b(new_n47_), .O(new_n218_));
  AND      g0202(.a(new_n83_), .b(i_2_3_99_0), .O(new_n219_));
  OR       g0203(.a(new_n219_), .b(new_n213_), .O(new_n220_));
  OR       g0204(.a(new_n220_), .b(new_n218_), .O(new_n221_));
  AND      g0205(.a(new_n221_), .b(new_n20_), .O(new_n222_));
  NOT      g0206(.a(i_2_3_68_0), .O(new_n223_));
  AND      g0207(.a(new_n223_), .b(i_2_3_43_0), .O(new_n224_));
  OR       g0208(.a(new_n132_), .b(i_2_3_42_0), .O(new_n225_));
  OR       g0209(.a(new_n225_), .b(i_2_3_79_0), .O(new_n226_));
  NAND     g0210(.a(new_n226_), .b(new_n101_), .O(new_n227_));
  AND      g0211(.a(new_n227_), .b(new_n224_), .O(new_n228_));
  OR       g0212(.a(new_n41_), .b(i_2_3_55_0), .O(new_n229_));
  NOT      g0213(.a(new_n96_), .O(new_n230_));
  AND      g0214(.a(new_n230_), .b(i_2_3_72_0), .O(new_n231_));
  AND      g0215(.a(new_n231_), .b(new_n229_), .O(new_n232_));
  OR       g0216(.a(new_n232_), .b(new_n228_), .O(new_n233_));
  OR       g0217(.a(new_n233_), .b(new_n222_), .O(new_n234_));
  AND      g0218(.a(new_n234_), .b(i_2_3_91_0), .O(new_n235_));
  AND      g0219(.a(new_n206_), .b(new_n53_), .O(new_n236_));
  OR       g0220(.a(i_2_3_72_0), .b(new_n77_), .O(new_n237_));
  OR       g0221(.a(new_n237_), .b(new_n212_), .O(new_n238_));
  AND      g0222(.a(new_n238_), .b(new_n236_), .O(new_n239_));
  OR       g0223(.a(new_n239_), .b(new_n219_), .O(new_n240_));
  AND      g0224(.a(new_n240_), .b(i_2_3_86_0), .O(new_n241_));
  OR       g0225(.a(new_n236_), .b(i_2_3_86_0), .O(new_n242_));
  AND      g0226(.a(new_n242_), .b(new_n31_), .O(new_n243_));
  OR       g0227(.a(new_n212_), .b(new_n31_), .O(new_n244_));
  NOT      g0228(.a(new_n34_), .O(new_n245_));
  AND      g0229(.a(new_n245_), .b(i_2_3_72_0), .O(new_n246_));
  AND      g0230(.a(new_n246_), .b(new_n244_), .O(new_n247_));
  OR       g0231(.a(new_n247_), .b(new_n243_), .O(new_n248_));
  OR       g0232(.a(new_n248_), .b(new_n241_), .O(new_n249_));
  AND      g0233(.a(new_n249_), .b(i_2_3_55_0), .O(new_n250_));
  OR       g0234(.a(i_2_3_55_0), .b(new_n53_), .O(new_n251_));
  NAND     g0235(.a(new_n251_), .b(new_n219_), .O(new_n252_));
  OR       g0236(.a(i_2_3_99_0), .b(i_2_3_43_0), .O(new_n253_));
  NAND     g0237(.a(new_n253_), .b(new_n237_), .O(new_n254_));
  AND      g0238(.a(new_n254_), .b(i_2_3_42_0), .O(new_n255_));
  NAND     g0239(.a(new_n237_), .b(new_n42_), .O(new_n256_));
  NAND     g0240(.a(new_n256_), .b(i_2_3_86_0), .O(new_n257_));
  OR       g0241(.a(new_n257_), .b(new_n255_), .O(new_n258_));
  NAND     g0242(.a(new_n258_), .b(new_n252_), .O(new_n259_));
  AND      g0243(.a(new_n259_), .b(new_n31_), .O(new_n260_));
  OR       g0244(.a(new_n260_), .b(new_n250_), .O(new_n261_));
  AND      g0245(.a(new_n261_), .b(new_n20_), .O(new_n262_));
  OR       g0246(.a(new_n262_), .b(new_n235_), .O(new_n263_));
  OR       g0247(.a(new_n263_), .b(new_n217_), .O(new_n264_));
  AND      g0248(.a(new_n264_), .b(i_2_3_29_0), .O(new_n265_));
  OR       g0249(.a(i_2_3_138_0), .b(i_2_3_43_0), .O(new_n266_));
  NOT      g0250(.a(new_n266_), .O(new_n267_));
  AND      g0251(.a(i_2_3_91_0), .b(i_2_3_43_0), .O(new_n268_));
  OR       g0252(.a(new_n268_), .b(new_n267_), .O(new_n269_));
  AND      g0253(.a(new_n269_), .b(i_2_3_55_0), .O(new_n270_));
  OR       g0254(.a(new_n270_), .b(new_n154_), .O(new_n271_));
  AND      g0255(.a(new_n271_), .b(new_n53_), .O(new_n272_));
  AND      g0256(.a(new_n200_), .b(new_n78_), .O(new_n273_));
  OR       g0257(.a(new_n273_), .b(new_n272_), .O(new_n274_));
  AND      g0258(.a(new_n274_), .b(new_n31_), .O(new_n275_));
  NAND     g0259(.a(new_n121_), .b(i_2_3_55_0), .O(new_n276_));
  AND      g0260(.a(new_n276_), .b(i_2_3_42_0), .O(new_n277_));
  OR       g0261(.a(i_2_3_79_0), .b(i_2_3_68_0), .O(new_n278_));
  OR       g0262(.a(new_n31_), .b(i_2_3_29_0), .O(new_n279_));
  OR       g0263(.a(new_n279_), .b(new_n278_), .O(new_n280_));
  AND      g0264(.a(new_n280_), .b(new_n132_), .O(new_n281_));
  OR       g0265(.a(new_n281_), .b(new_n24_), .O(new_n282_));
  OR       g0266(.a(new_n282_), .b(new_n277_), .O(new_n283_));
  OR       g0267(.a(new_n278_), .b(i_2_3_138_0), .O(new_n284_));
  OR       g0268(.a(new_n284_), .b(new_n23_), .O(new_n285_));
  NAND     g0269(.a(new_n285_), .b(new_n283_), .O(new_n286_));
  AND      g0270(.a(new_n286_), .b(i_2_3_99_0), .O(new_n287_));
  OR       g0271(.a(new_n287_), .b(new_n275_), .O(new_n288_));
  AND      g0272(.a(new_n288_), .b(i_2_3_72_0), .O(new_n289_));
  AND      g0273(.a(new_n67_), .b(new_n206_), .O(new_n290_));
  OR       g0274(.a(new_n268_), .b(new_n256_), .O(new_n291_));
  AND      g0275(.a(new_n71_), .b(new_n31_), .O(new_n292_));
  AND      g0276(.a(new_n292_), .b(new_n291_), .O(new_n293_));
  OR       g0277(.a(new_n293_), .b(new_n290_), .O(new_n294_));
  AND      g0278(.a(new_n294_), .b(new_n20_), .O(new_n295_));
  AND      g0279(.a(new_n213_), .b(new_n76_), .O(new_n296_));
  OR       g0280(.a(new_n296_), .b(new_n295_), .O(new_n297_));
  AND      g0281(.a(new_n297_), .b(new_n53_), .O(new_n298_));
  OR       g0282(.a(new_n298_), .b(new_n289_), .O(new_n299_));
  AND      g0283(.a(new_n299_), .b(i_2_3_86_0), .O(new_n300_));
  AND      g0284(.a(new_n20_), .b(i_2_3_43_0), .O(new_n301_));
  AND      g0285(.a(new_n301_), .b(new_n129_), .O(new_n302_));
  OR       g0286(.a(i_2_3_99_0), .b(i_2_3_72_0), .O(new_n303_));
  AND      g0287(.a(new_n303_), .b(new_n154_), .O(new_n304_));
  AND      g0288(.a(new_n20_), .b(i_2_3_99_0), .O(new_n305_));
  AND      g0289(.a(new_n78_), .b(new_n40_), .O(new_n306_));
  OR       g0290(.a(new_n306_), .b(new_n305_), .O(new_n307_));
  AND      g0291(.a(new_n307_), .b(new_n83_), .O(new_n308_));
  OR       g0292(.a(new_n308_), .b(new_n304_), .O(new_n309_));
  AND      g0293(.a(new_n309_), .b(new_n53_), .O(new_n310_));
  OR       g0294(.a(i_2_3_79_0), .b(i_2_3_72_0), .O(new_n311_));
  NOT      g0295(.a(new_n311_), .O(new_n312_));
  AND      g0296(.a(new_n312_), .b(new_n154_), .O(new_n313_));
  OR       g0297(.a(new_n313_), .b(new_n310_), .O(new_n314_));
  AND      g0298(.a(new_n314_), .b(i_2_3_55_0), .O(new_n315_));
  AND      g0299(.a(new_n83_), .b(new_n20_), .O(new_n316_));
  AND      g0300(.a(i_2_3_99_0), .b(i_2_3_91_0), .O(new_n317_));
  AND      g0301(.a(new_n317_), .b(new_n316_), .O(new_n318_));
  OR       g0302(.a(new_n318_), .b(new_n315_), .O(new_n319_));
  AND      g0303(.a(new_n319_), .b(new_n31_), .O(new_n320_));
  OR       g0304(.a(new_n320_), .b(new_n302_), .O(new_n321_));
  OR       g0305(.a(new_n321_), .b(new_n300_), .O(new_n322_));
  OR       g0306(.a(new_n322_), .b(new_n265_), .O(new_n323_));
  OR       g0307(.a(new_n323_), .b(new_n191_), .O(new_n324_));
  AND      g0308(.a(new_n324_), .b(new_n19_), .O(new_n325_));
  AND      g0309(.a(i_2_3_86_0), .b(new_n53_), .O(new_n326_));
  AND      g0310(.a(new_n200_), .b(i_2_3_99_0), .O(new_n327_));
  OR       g0311(.a(new_n327_), .b(new_n326_), .O(new_n328_));
  AND      g0312(.a(new_n328_), .b(new_n56_), .O(new_n329_));
  NOT      g0313(.a(new_n225_), .O(new_n330_));
  AND      g0314(.a(new_n22_), .b(i_2_3_29_0), .O(new_n331_));
  OR       g0315(.a(new_n331_), .b(new_n330_), .O(new_n332_));
  NAND     g0316(.a(new_n332_), .b(new_n31_), .O(new_n333_));
  NAND     g0317(.a(i_2_3_99_0), .b(i_2_3_77_0), .O(new_n334_));
  OR       g0318(.a(new_n334_), .b(new_n69_), .O(new_n335_));
  NAND     g0319(.a(new_n335_), .b(new_n333_), .O(new_n336_));
  OR       g0320(.a(new_n336_), .b(new_n329_), .O(new_n337_));
  AND      g0321(.a(new_n337_), .b(i_2_3_72_0), .O(new_n338_));
  AND      g0322(.a(new_n326_), .b(new_n147_), .O(new_n339_));
  AND      g0323(.a(new_n99_), .b(i_2_3_72_0), .O(new_n340_));
  NOT      g0324(.a(new_n340_), .O(new_n341_));
  AND      g0325(.a(new_n303_), .b(i_2_3_55_0), .O(new_n342_));
  AND      g0326(.a(new_n342_), .b(new_n341_), .O(new_n343_));
  OR       g0327(.a(new_n343_), .b(new_n339_), .O(new_n344_));
  AND      g0328(.a(new_n344_), .b(new_n279_), .O(new_n345_));
  OR       g0329(.a(new_n226_), .b(new_n99_), .O(new_n346_));
  AND      g0330(.a(new_n200_), .b(i_2_3_86_0), .O(new_n347_));
  AND      g0331(.a(i_2_3_99_0), .b(new_n53_), .O(new_n348_));
  OR       g0332(.a(new_n348_), .b(new_n347_), .O(new_n349_));
  NAND     g0333(.a(new_n349_), .b(i_2_3_29_0), .O(new_n350_));
  NAND     g0334(.a(new_n350_), .b(new_n346_), .O(new_n351_));
  AND      g0335(.a(new_n128_), .b(i_2_3_86_0), .O(new_n352_));
  AND      g0336(.a(i_2_3_99_0), .b(new_n31_), .O(new_n353_));
  OR       g0337(.a(new_n353_), .b(new_n352_), .O(new_n354_));
  AND      g0338(.a(i_2_3_99_0), .b(i_2_3_86_0), .O(new_n355_));
  NOT      g0339(.a(new_n355_), .O(new_n356_));
  AND      g0340(.a(new_n356_), .b(i_2_3_43_0), .O(new_n357_));
  AND      g0341(.a(new_n357_), .b(new_n354_), .O(new_n358_));
  NOT      g0342(.a(i_2_3_29_0), .O(new_n359_));
  AND      g0343(.a(new_n356_), .b(new_n359_), .O(new_n360_));
  NAND     g0344(.a(new_n360_), .b(new_n226_), .O(new_n361_));
  AND      g0345(.a(new_n63_), .b(new_n31_), .O(new_n362_));
  AND      g0346(.a(new_n362_), .b(new_n361_), .O(new_n363_));
  OR       g0347(.a(new_n363_), .b(new_n358_), .O(new_n364_));
  OR       g0348(.a(new_n364_), .b(new_n351_), .O(new_n365_));
  OR       g0349(.a(new_n365_), .b(new_n345_), .O(new_n366_));
  OR       g0350(.a(new_n366_), .b(new_n338_), .O(new_n367_));
  AND      g0351(.a(new_n367_), .b(i_2_3_68_0), .O(new_n368_));
  AND      g0352(.a(new_n19_), .b(i_2_3_72_0), .O(new_n369_));
  NOT      g0353(.a(new_n369_), .O(new_n370_));
  OR       g0354(.a(new_n166_), .b(i_2_3_72_0), .O(new_n371_));
  NAND     g0355(.a(new_n371_), .b(i_2_3_79_0), .O(new_n372_));
  AND      g0356(.a(new_n372_), .b(new_n370_), .O(new_n373_));
  AND      g0357(.a(i_2_3_99_0), .b(i_2_3_72_0), .O(new_n374_));
  OR       g0358(.a(new_n374_), .b(new_n54_), .O(new_n375_));
  OR       g0359(.a(new_n375_), .b(new_n373_), .O(new_n376_));
  AND      g0360(.a(new_n376_), .b(i_2_3_29_0), .O(new_n377_));
  AND      g0361(.a(new_n206_), .b(i_2_3_86_0), .O(new_n378_));
  NAND     g0362(.a(new_n34_), .b(new_n132_), .O(new_n379_));
  AND      g0363(.a(new_n379_), .b(new_n378_), .O(new_n380_));
  AND      g0364(.a(i_2_3_99_0), .b(new_n77_), .O(new_n381_));
  OR       g0365(.a(new_n381_), .b(new_n21_), .O(new_n382_));
  AND      g0366(.a(new_n382_), .b(new_n330_), .O(new_n383_));
  OR       g0367(.a(new_n383_), .b(new_n380_), .O(new_n384_));
  AND      g0368(.a(new_n384_), .b(i_2_3_72_0), .O(new_n385_));
  OR       g0369(.a(new_n212_), .b(i_2_3_55_0), .O(new_n386_));
  AND      g0370(.a(new_n386_), .b(new_n328_), .O(new_n387_));
  OR       g0371(.a(new_n387_), .b(new_n385_), .O(new_n388_));
  OR       g0372(.a(new_n388_), .b(new_n377_), .O(new_n389_));
  AND      g0373(.a(new_n389_), .b(new_n31_), .O(new_n390_));
  OR       g0374(.a(new_n178_), .b(i_2_3_72_0), .O(new_n391_));
  AND      g0375(.a(new_n348_), .b(new_n200_), .O(new_n392_));
  AND      g0376(.a(new_n392_), .b(new_n391_), .O(new_n393_));
  OR       g0377(.a(new_n374_), .b(new_n56_), .O(new_n394_));
  AND      g0378(.a(new_n394_), .b(new_n77_), .O(new_n395_));
  OR       g0379(.a(new_n56_), .b(i_2_3_77_0), .O(new_n396_));
  AND      g0380(.a(new_n396_), .b(new_n395_), .O(new_n397_));
  AND      g0381(.a(new_n56_), .b(i_2_3_99_0), .O(new_n398_));
  OR       g0382(.a(new_n398_), .b(new_n139_), .O(new_n399_));
  OR       g0383(.a(i_2_3_99_0), .b(i_2_3_86_0), .O(new_n400_));
  OR       g0384(.a(new_n355_), .b(i_2_3_55_0), .O(new_n401_));
  AND      g0385(.a(new_n401_), .b(new_n400_), .O(new_n402_));
  AND      g0386(.a(new_n402_), .b(new_n399_), .O(new_n403_));
  OR       g0387(.a(new_n403_), .b(new_n397_), .O(new_n404_));
  AND      g0388(.a(new_n404_), .b(new_n53_), .O(new_n405_));
  NOT      g0389(.a(new_n100_), .O(new_n406_));
  AND      g0390(.a(new_n342_), .b(new_n406_), .O(new_n407_));
  OR       g0391(.a(new_n407_), .b(new_n405_), .O(new_n408_));
  AND      g0392(.a(new_n408_), .b(i_2_3_29_0), .O(new_n409_));
  OR       g0393(.a(new_n409_), .b(new_n393_), .O(new_n410_));
  OR       g0394(.a(new_n410_), .b(new_n390_), .O(new_n411_));
  OR       g0395(.a(new_n411_), .b(new_n368_), .O(new_n412_));
  AND      g0396(.a(new_n412_), .b(i_2_3_91_0), .O(new_n413_));
  NOT      g0397(.a(new_n56_), .O(new_n414_));
  NAND     g0398(.a(new_n225_), .b(new_n414_), .O(new_n415_));
  OR       g0399(.a(new_n326_), .b(i_2_3_29_0), .O(new_n416_));
  AND      g0400(.a(new_n416_), .b(new_n415_), .O(new_n417_));
  OR       g0401(.a(new_n56_), .b(new_n54_), .O(new_n418_));
  AND      g0402(.a(new_n418_), .b(i_2_3_72_0), .O(new_n419_));
  OR       g0403(.a(i_2_3_86_0), .b(new_n132_), .O(new_n420_));
  AND      g0404(.a(new_n420_), .b(i_2_3_43_0), .O(new_n421_));
  OR       g0405(.a(new_n421_), .b(new_n183_), .O(new_n422_));
  OR       g0406(.a(new_n422_), .b(new_n419_), .O(new_n423_));
  AND      g0407(.a(new_n423_), .b(i_2_3_99_0), .O(new_n424_));
  OR       g0408(.a(new_n424_), .b(new_n417_), .O(new_n425_));
  AND      g0409(.a(new_n425_), .b(new_n21_), .O(new_n426_));
  AND      g0410(.a(new_n30_), .b(i_2_3_86_0), .O(new_n427_));
  AND      g0411(.a(new_n427_), .b(i_2_3_29_0), .O(new_n428_));
  AND      g0412(.a(new_n331_), .b(new_n303_), .O(new_n429_));
  AND      g0413(.a(i_2_3_72_0), .b(new_n77_), .O(new_n430_));
  OR       g0414(.a(new_n430_), .b(i_2_3_99_0), .O(new_n431_));
  AND      g0415(.a(new_n431_), .b(new_n56_), .O(new_n432_));
  OR       g0416(.a(new_n432_), .b(new_n429_), .O(new_n433_));
  AND      g0417(.a(new_n433_), .b(new_n53_), .O(new_n434_));
  OR       g0418(.a(new_n434_), .b(new_n428_), .O(new_n435_));
  OR       g0419(.a(new_n435_), .b(new_n426_), .O(new_n436_));
  AND      g0420(.a(new_n436_), .b(i_2_3_68_0), .O(new_n437_));
  AND      g0421(.a(new_n393_), .b(i_2_3_86_0), .O(new_n438_));
  OR       g0422(.a(new_n278_), .b(new_n99_), .O(new_n439_));
  OR       g0423(.a(new_n225_), .b(new_n25_), .O(new_n440_));
  NAND     g0424(.a(new_n440_), .b(new_n439_), .O(new_n441_));
  AND      g0425(.a(new_n441_), .b(i_2_3_99_0), .O(new_n442_));
  OR       g0426(.a(new_n326_), .b(new_n83_), .O(new_n443_));
  AND      g0427(.a(new_n443_), .b(new_n415_), .O(new_n444_));
  OR       g0428(.a(new_n444_), .b(new_n442_), .O(new_n445_));
  AND      g0429(.a(new_n445_), .b(new_n77_), .O(new_n446_));
  AND      g0430(.a(new_n303_), .b(new_n330_), .O(new_n447_));
  OR       g0431(.a(new_n447_), .b(new_n219_), .O(new_n448_));
  AND      g0432(.a(new_n448_), .b(i_2_3_86_0), .O(new_n449_));
  OR       g0433(.a(new_n449_), .b(new_n392_), .O(new_n450_));
  OR       g0434(.a(new_n450_), .b(new_n446_), .O(new_n451_));
  AND      g0435(.a(new_n451_), .b(i_2_3_29_0), .O(new_n452_));
  OR       g0436(.a(new_n452_), .b(new_n438_), .O(new_n453_));
  OR       g0437(.a(new_n453_), .b(new_n437_), .O(new_n454_));
  AND      g0438(.a(new_n454_), .b(new_n31_), .O(new_n455_));
  OR       g0439(.a(new_n34_), .b(new_n132_), .O(new_n456_));
  NAND     g0440(.a(new_n456_), .b(new_n359_), .O(new_n457_));
  AND      g0441(.a(i_2_3_99_0), .b(i_2_3_68_0), .O(new_n458_));
  AND      g0442(.a(new_n458_), .b(i_2_3_72_0), .O(new_n459_));
  AND      g0443(.a(new_n459_), .b(new_n406_), .O(new_n460_));
  AND      g0444(.a(new_n460_), .b(new_n457_), .O(new_n461_));
  AND      g0445(.a(new_n458_), .b(new_n83_), .O(new_n462_));
  NOT      g0446(.a(new_n219_), .O(new_n463_));
  AND      g0447(.a(new_n206_), .b(i_2_3_68_0), .O(new_n464_));
  NOT      g0448(.a(new_n464_), .O(new_n465_));
  AND      g0449(.a(new_n465_), .b(new_n463_), .O(new_n466_));
  OR       g0450(.a(new_n430_), .b(new_n212_), .O(new_n467_));
  OR       g0451(.a(new_n212_), .b(i_2_3_68_0), .O(new_n468_));
  AND      g0452(.a(new_n468_), .b(new_n77_), .O(new_n469_));
  NAND     g0453(.a(new_n469_), .b(new_n467_), .O(new_n470_));
  NAND     g0454(.a(new_n470_), .b(new_n466_), .O(new_n471_));
  AND      g0455(.a(new_n471_), .b(i_2_3_86_0), .O(new_n472_));
  OR       g0456(.a(new_n472_), .b(new_n462_), .O(new_n473_));
  AND      g0457(.a(new_n330_), .b(i_2_3_29_0), .O(new_n474_));
  AND      g0458(.a(new_n474_), .b(new_n473_), .O(new_n475_));
  OR       g0459(.a(new_n475_), .b(new_n461_), .O(new_n476_));
  OR       g0460(.a(new_n476_), .b(new_n455_), .O(new_n477_));
  OR       g0461(.a(new_n477_), .b(new_n413_), .O(new_n478_));
  AND      g0462(.a(new_n478_), .b(new_n20_), .O(new_n479_));
  OR       g0463(.a(new_n25_), .b(i_2_3_43_0), .O(new_n480_));
  OR       g0464(.a(new_n480_), .b(i_2_3_68_0), .O(new_n481_));
  AND      g0465(.a(new_n481_), .b(new_n398_), .O(new_n482_));
  AND      g0466(.a(new_n25_), .b(i_2_3_68_0), .O(new_n483_));
  AND      g0467(.a(new_n483_), .b(i_2_3_99_0), .O(new_n484_));
  OR       g0468(.a(new_n484_), .b(new_n427_), .O(new_n485_));
  OR       g0469(.a(new_n485_), .b(new_n397_), .O(new_n486_));
  AND      g0470(.a(new_n486_), .b(new_n21_), .O(new_n487_));
  OR       g0471(.a(new_n487_), .b(new_n482_), .O(new_n488_));
  AND      g0472(.a(new_n488_), .b(new_n31_), .O(new_n489_));
  AND      g0473(.a(new_n402_), .b(new_n31_), .O(new_n490_));
  AND      g0474(.a(new_n398_), .b(i_2_3_72_0), .O(new_n491_));
  OR       g0475(.a(new_n491_), .b(new_n490_), .O(new_n492_));
  AND      g0476(.a(new_n492_), .b(i_2_3_68_0), .O(new_n493_));
  OR       g0477(.a(new_n109_), .b(i_2_3_72_0), .O(new_n494_));
  AND      g0478(.a(new_n494_), .b(i_2_3_43_0), .O(new_n495_));
  AND      g0479(.a(new_n483_), .b(i_2_3_55_0), .O(new_n496_));
  OR       g0480(.a(new_n496_), .b(new_n495_), .O(new_n497_));
  AND      g0481(.a(new_n497_), .b(i_2_3_99_0), .O(new_n498_));
  AND      g0482(.a(i_2_3_68_0), .b(new_n31_), .O(new_n499_));
  AND      g0483(.a(new_n22_), .b(new_n77_), .O(new_n500_));
  OR       g0484(.a(new_n500_), .b(new_n66_), .O(new_n501_));
  AND      g0485(.a(new_n501_), .b(new_n499_), .O(new_n502_));
  OR       g0486(.a(new_n502_), .b(new_n427_), .O(new_n503_));
  OR       g0487(.a(new_n503_), .b(new_n498_), .O(new_n504_));
  AND      g0488(.a(new_n504_), .b(new_n21_), .O(new_n505_));
  OR       g0489(.a(new_n505_), .b(new_n493_), .O(new_n506_));
  AND      g0490(.a(new_n506_), .b(new_n53_), .O(new_n507_));
  OR       g0491(.a(new_n507_), .b(new_n489_), .O(new_n508_));
  AND      g0492(.a(new_n508_), .b(i_2_3_91_0), .O(new_n509_));
  NOT      g0493(.a(new_n458_), .O(new_n510_));
  AND      g0494(.a(new_n21_), .b(i_2_3_68_0), .O(new_n511_));
  NAND     g0495(.a(new_n511_), .b(i_2_3_72_0), .O(new_n512_));
  NAND     g0496(.a(new_n512_), .b(new_n510_), .O(new_n513_));
  AND      g0497(.a(new_n339_), .b(new_n213_), .O(new_n514_));
  AND      g0498(.a(new_n514_), .b(new_n513_), .O(new_n515_));
  OR       g0499(.a(new_n515_), .b(new_n509_), .O(new_n516_));
  AND      g0500(.a(new_n516_), .b(i_2_3_29_0), .O(new_n517_));
  NOT      g0501(.a(new_n466_), .O(new_n518_));
  AND      g0502(.a(new_n518_), .b(new_n52_), .O(new_n519_));
  AND      g0503(.a(new_n519_), .b(new_n329_), .O(new_n520_));
  OR       g0504(.a(new_n520_), .b(new_n517_), .O(new_n521_));
  OR       g0505(.a(new_n521_), .b(new_n479_), .O(new_n522_));
  OR       g0506(.a(new_n522_), .b(new_n325_), .O(new_n523_));
  AND      g0507(.a(new_n523_), .b(new_n18_), .O(new_n524_));
  AND      g0508(.a(i_2_3_99_0), .b(new_n19_), .O(new_n525_));
  OR       g0509(.a(new_n525_), .b(new_n31_), .O(new_n526_));
  AND      g0510(.a(new_n526_), .b(i_2_3_55_0), .O(new_n527_));
  AND      g0511(.a(i_2_3_143_0), .b(new_n77_), .O(new_n528_));
  AND      g0512(.a(new_n528_), .b(i_2_3_68_0), .O(new_n529_));
  OR       g0513(.a(new_n529_), .b(new_n78_), .O(new_n530_));
  OR       g0514(.a(new_n530_), .b(new_n527_), .O(new_n531_));
  AND      g0515(.a(new_n531_), .b(i_2_3_86_0), .O(new_n532_));
  AND      g0516(.a(new_n19_), .b(i_2_3_68_0), .O(new_n533_));
  AND      g0517(.a(new_n533_), .b(i_2_3_143_0), .O(new_n534_));
  AND      g0518(.a(new_n534_), .b(i_2_3_99_0), .O(new_n535_));
  OR       g0519(.a(new_n535_), .b(new_n67_), .O(new_n536_));
  OR       g0520(.a(new_n536_), .b(new_n532_), .O(new_n537_));
  AND      g0521(.a(new_n537_), .b(new_n20_), .O(new_n538_));
  AND      g0522(.a(i_2_3_143_0), .b(new_n19_), .O(new_n539_));
  AND      g0523(.a(new_n178_), .b(new_n20_), .O(new_n540_));
  NAND     g0524(.a(new_n540_), .b(new_n539_), .O(new_n541_));
  OR       g0525(.a(new_n400_), .b(i_2_3_68_0), .O(new_n542_));
  OR       g0526(.a(new_n542_), .b(new_n118_), .O(new_n543_));
  NAND     g0527(.a(new_n543_), .b(new_n541_), .O(new_n544_));
  AND      g0528(.a(new_n544_), .b(new_n132_), .O(new_n545_));
  NAND     g0529(.a(i_2_3_143_0), .b(i_2_3_77_0), .O(new_n546_));
  NOT      g0530(.a(new_n546_), .O(new_n547_));
  AND      g0531(.a(new_n547_), .b(new_n317_), .O(new_n548_));
  OR       g0532(.a(i_2_3_99_0), .b(new_n19_), .O(new_n549_));
  AND      g0533(.a(new_n549_), .b(i_2_3_55_0), .O(new_n550_));
  AND      g0534(.a(new_n550_), .b(new_n31_), .O(new_n551_));
  OR       g0535(.a(new_n551_), .b(new_n548_), .O(new_n552_));
  AND      g0536(.a(new_n552_), .b(i_2_3_68_0), .O(new_n553_));
  AND      g0537(.a(new_n224_), .b(i_2_3_138_0), .O(new_n554_));
  OR       g0538(.a(new_n499_), .b(i_2_3_55_0), .O(new_n555_));
  OR       g0539(.a(new_n555_), .b(new_n554_), .O(new_n556_));
  AND      g0540(.a(i_2_3_91_0), .b(new_n19_), .O(new_n557_));
  AND      g0541(.a(new_n557_), .b(new_n556_), .O(new_n558_));
  OR       g0542(.a(new_n558_), .b(new_n553_), .O(new_n559_));
  AND      g0543(.a(new_n559_), .b(i_2_3_86_0), .O(new_n560_));
  OR       g0544(.a(new_n560_), .b(new_n545_), .O(new_n561_));
  OR       g0545(.a(new_n561_), .b(new_n538_), .O(new_n562_));
  AND      g0546(.a(new_n562_), .b(new_n21_), .O(new_n563_));
  AND      g0547(.a(i_2_3_68_0), .b(i_2_3_55_0), .O(new_n564_));
  AND      g0548(.a(new_n564_), .b(new_n20_), .O(new_n565_));
  AND      g0549(.a(new_n20_), .b(i_2_3_55_0), .O(new_n566_));
  AND      g0550(.a(new_n317_), .b(i_2_3_68_0), .O(new_n567_));
  OR       g0551(.a(new_n567_), .b(new_n566_), .O(new_n568_));
  AND      g0552(.a(new_n568_), .b(new_n77_), .O(new_n569_));
  AND      g0553(.a(new_n317_), .b(i_2_3_55_0), .O(new_n570_));
  OR       g0554(.a(new_n570_), .b(new_n569_), .O(new_n571_));
  AND      g0555(.a(new_n571_), .b(new_n19_), .O(new_n572_));
  OR       g0556(.a(new_n572_), .b(new_n565_), .O(new_n573_));
  AND      g0557(.a(new_n573_), .b(new_n21_), .O(new_n574_));
  AND      g0558(.a(i_2_3_86_0), .b(new_n19_), .O(new_n575_));
  AND      g0559(.a(new_n575_), .b(new_n567_), .O(new_n576_));
  AND      g0560(.a(i_2_3_86_0), .b(i_2_3_68_0), .O(new_n577_));
  OR       g0561(.a(new_n525_), .b(i_2_3_91_0), .O(new_n578_));
  AND      g0562(.a(new_n578_), .b(new_n577_), .O(new_n579_));
  OR       g0563(.a(new_n533_), .b(new_n355_), .O(new_n580_));
  AND      g0564(.a(new_n580_), .b(new_n78_), .O(new_n581_));
  OR       g0565(.a(new_n581_), .b(new_n579_), .O(new_n582_));
  AND      g0566(.a(new_n582_), .b(i_2_3_55_0), .O(new_n583_));
  OR       g0567(.a(new_n583_), .b(new_n576_), .O(new_n584_));
  OR       g0568(.a(new_n584_), .b(new_n574_), .O(new_n585_));
  AND      g0569(.a(new_n585_), .b(new_n31_), .O(new_n586_));
  NAND     g0570(.a(i_2_3_143_0), .b(i_2_3_99_0), .O(new_n587_));
  NAND     g0571(.a(new_n587_), .b(i_2_3_77_0), .O(new_n588_));
  OR       g0572(.a(new_n588_), .b(i_2_3_68_0), .O(new_n589_));
  AND      g0573(.a(new_n589_), .b(i_2_3_55_0), .O(new_n590_));
  OR       g0574(.a(new_n42_), .b(new_n77_), .O(new_n591_));
  AND      g0575(.a(new_n591_), .b(new_n575_), .O(new_n592_));
  OR       g0576(.a(new_n592_), .b(new_n534_), .O(new_n593_));
  OR       g0577(.a(new_n593_), .b(new_n590_), .O(new_n594_));
  AND      g0578(.a(new_n594_), .b(i_2_3_91_0), .O(new_n595_));
  NOT      g0579(.a(new_n575_), .O(new_n596_));
  OR       g0580(.a(new_n18_), .b(i_2_3_43_0), .O(new_n597_));
  OR       g0581(.a(new_n597_), .b(new_n334_), .O(new_n598_));
  NAND     g0582(.a(new_n598_), .b(new_n596_), .O(new_n599_));
  AND      g0583(.a(new_n599_), .b(new_n31_), .O(new_n600_));
  OR       g0584(.a(new_n213_), .b(new_n178_), .O(new_n601_));
  AND      g0585(.a(new_n601_), .b(new_n550_), .O(new_n602_));
  OR       g0586(.a(new_n602_), .b(new_n600_), .O(new_n603_));
  AND      g0587(.a(new_n603_), .b(i_2_3_68_0), .O(new_n604_));
  AND      g0588(.a(new_n578_), .b(new_n500_), .O(new_n605_));
  AND      g0589(.a(new_n550_), .b(i_2_3_86_0), .O(new_n606_));
  OR       g0590(.a(new_n606_), .b(new_n605_), .O(new_n607_));
  AND      g0591(.a(new_n607_), .b(new_n31_), .O(new_n608_));
  OR       g0592(.a(new_n608_), .b(new_n604_), .O(new_n609_));
  OR       g0593(.a(new_n609_), .b(new_n595_), .O(new_n610_));
  AND      g0594(.a(new_n610_), .b(new_n20_), .O(new_n611_));
  OR       g0595(.a(new_n611_), .b(new_n586_), .O(new_n612_));
  OR       g0596(.a(new_n612_), .b(new_n563_), .O(new_n613_));
  AND      g0597(.a(new_n613_), .b(i_2_3_72_0), .O(new_n614_));
  OR       g0598(.a(new_n212_), .b(new_n77_), .O(new_n615_));
  AND      g0599(.a(new_n615_), .b(new_n378_), .O(new_n616_));
  AND      g0600(.a(new_n32_), .b(new_n19_), .O(new_n617_));
  OR       g0601(.a(new_n511_), .b(new_n353_), .O(new_n618_));
  OR       g0602(.a(new_n618_), .b(new_n577_), .O(new_n619_));
  OR       g0603(.a(new_n619_), .b(new_n617_), .O(new_n620_));
  OR       g0604(.a(new_n620_), .b(new_n616_), .O(new_n621_));
  AND      g0605(.a(new_n621_), .b(i_2_3_91_0), .O(new_n622_));
  AND      g0606(.a(new_n244_), .b(i_2_3_68_0), .O(new_n623_));
  NAND     g0607(.a(i_2_3_79_0), .b(i_2_3_77_0), .O(new_n624_));
  AND      g0608(.a(new_n624_), .b(i_2_3_99_0), .O(new_n625_));
  OR       g0609(.a(i_2_3_77_0), .b(i_2_3_43_0), .O(new_n626_));
  OR       g0610(.a(new_n626_), .b(i_2_3_79_0), .O(new_n627_));
  NAND     g0611(.a(new_n627_), .b(i_2_3_47_0), .O(new_n628_));
  AND      g0612(.a(new_n628_), .b(new_n625_), .O(new_n629_));
  OR       g0613(.a(new_n629_), .b(new_n623_), .O(new_n630_));
  AND      g0614(.a(new_n630_), .b(i_2_3_86_0), .O(new_n631_));
  OR       g0615(.a(i_2_3_79_0), .b(i_2_3_77_0), .O(new_n632_));
  NOT      g0616(.a(new_n632_), .O(new_n633_));
  AND      g0617(.a(new_n633_), .b(new_n353_), .O(new_n634_));
  OR       g0618(.a(new_n533_), .b(new_n179_), .O(new_n635_));
  AND      g0619(.a(new_n206_), .b(new_n32_), .O(new_n636_));
  AND      g0620(.a(new_n636_), .b(new_n635_), .O(new_n637_));
  OR       g0621(.a(new_n637_), .b(new_n634_), .O(new_n638_));
  OR       g0622(.a(new_n638_), .b(new_n631_), .O(new_n639_));
  OR       g0623(.a(new_n639_), .b(new_n622_), .O(new_n640_));
  AND      g0624(.a(new_n640_), .b(i_2_3_55_0), .O(new_n641_));
  OR       g0625(.a(new_n21_), .b(i_2_3_68_0), .O(new_n642_));
  AND      g0626(.a(new_n642_), .b(new_n525_), .O(new_n643_));
  AND      g0627(.a(new_n312_), .b(i_2_3_68_0), .O(new_n644_));
  OR       g0628(.a(new_n644_), .b(new_n643_), .O(new_n645_));
  AND      g0629(.a(new_n645_), .b(i_2_3_86_0), .O(new_n646_));
  AND      g0630(.a(new_n511_), .b(i_2_3_99_0), .O(new_n647_));
  AND      g0631(.a(new_n647_), .b(new_n547_), .O(new_n648_));
  OR       g0632(.a(new_n648_), .b(new_n646_), .O(new_n649_));
  AND      g0633(.a(new_n649_), .b(new_n31_), .O(new_n650_));
  NAND     g0634(.a(new_n632_), .b(new_n131_), .O(new_n651_));
  AND      g0635(.a(new_n651_), .b(new_n77_), .O(new_n652_));
  AND      g0636(.a(new_n525_), .b(i_2_3_86_0), .O(new_n653_));
  OR       g0637(.a(new_n653_), .b(new_n652_), .O(new_n654_));
  AND      g0638(.a(new_n654_), .b(i_2_3_68_0), .O(new_n655_));
  NAND     g0639(.a(new_n632_), .b(i_2_3_47_0), .O(new_n656_));
  AND      g0640(.a(new_n656_), .b(new_n355_), .O(new_n657_));
  AND      g0641(.a(new_n499_), .b(i_2_3_77_0), .O(new_n658_));
  AND      g0642(.a(new_n200_), .b(new_n99_), .O(new_n659_));
  OR       g0643(.a(new_n659_), .b(new_n658_), .O(new_n660_));
  AND      g0644(.a(new_n660_), .b(i_2_3_43_0), .O(new_n661_));
  OR       g0645(.a(new_n661_), .b(new_n657_), .O(new_n662_));
  OR       g0646(.a(new_n662_), .b(new_n655_), .O(new_n663_));
  AND      g0647(.a(new_n663_), .b(i_2_3_91_0), .O(new_n664_));
  OR       g0648(.a(new_n664_), .b(new_n650_), .O(new_n665_));
  OR       g0649(.a(new_n665_), .b(new_n641_), .O(new_n666_));
  AND      g0650(.a(new_n666_), .b(new_n20_), .O(new_n667_));
  AND      g0651(.a(new_n170_), .b(new_n19_), .O(new_n668_));
  AND      g0652(.a(new_n668_), .b(new_n601_), .O(new_n669_));
  OR       g0653(.a(new_n669_), .b(new_n214_), .O(new_n670_));
  AND      g0654(.a(new_n670_), .b(new_n206_), .O(new_n671_));
  AND      g0655(.a(new_n353_), .b(new_n139_), .O(new_n672_));
  OR       g0656(.a(new_n672_), .b(new_n671_), .O(new_n673_));
  AND      g0657(.a(new_n673_), .b(i_2_3_91_0), .O(new_n674_));
  AND      g0658(.a(new_n215_), .b(new_n19_), .O(new_n675_));
  OR       g0659(.a(new_n675_), .b(new_n674_), .O(new_n676_));
  AND      g0660(.a(new_n676_), .b(i_2_3_68_0), .O(new_n677_));
  AND      g0661(.a(new_n163_), .b(new_n19_), .O(new_n678_));
  OR       g0662(.a(new_n678_), .b(new_n677_), .O(new_n679_));
  OR       g0663(.a(new_n679_), .b(new_n667_), .O(new_n680_));
  OR       g0664(.a(new_n680_), .b(new_n614_), .O(new_n681_));
  AND      g0665(.a(new_n681_), .b(new_n53_), .O(new_n682_));
  AND      g0666(.a(new_n624_), .b(new_n56_), .O(new_n683_));
  NAND     g0667(.a(i_2_3_77_0), .b(i_2_3_55_0), .O(new_n684_));
  AND      g0668(.a(new_n684_), .b(new_n212_), .O(new_n685_));
  OR       g0669(.a(new_n685_), .b(new_n683_), .O(new_n686_));
  AND      g0670(.a(new_n686_), .b(i_2_3_68_0), .O(new_n687_));
  AND      g0671(.a(new_n19_), .b(i_2_3_55_0), .O(new_n688_));
  AND      g0672(.a(new_n688_), .b(new_n378_), .O(new_n689_));
  OR       g0673(.a(new_n689_), .b(new_n687_), .O(new_n690_));
  AND      g0674(.a(new_n690_), .b(i_2_3_72_0), .O(new_n691_));
  AND      g0675(.a(new_n615_), .b(new_n19_), .O(new_n692_));
  OR       g0676(.a(new_n692_), .b(new_n458_), .O(new_n693_));
  AND      g0677(.a(new_n693_), .b(new_n56_), .O(new_n694_));
  OR       g0678(.a(new_n694_), .b(new_n691_), .O(new_n695_));
  AND      g0679(.a(new_n695_), .b(new_n31_), .O(new_n696_));
  AND      g0680(.a(new_n193_), .b(i_2_3_99_0), .O(new_n697_));
  OR       g0681(.a(new_n549_), .b(i_2_3_79_0), .O(new_n698_));
  NAND     g0682(.a(new_n698_), .b(new_n356_), .O(new_n699_));
  AND      g0683(.a(new_n699_), .b(i_2_3_72_0), .O(new_n700_));
  OR       g0684(.a(new_n100_), .b(new_n40_), .O(new_n701_));
  NAND     g0685(.a(i_2_3_47_0), .b(i_2_3_43_0), .O(new_n702_));
  OR       g0686(.a(new_n702_), .b(new_n632_), .O(new_n703_));
  NAND     g0687(.a(new_n703_), .b(new_n701_), .O(new_n704_));
  OR       g0688(.a(new_n704_), .b(new_n700_), .O(new_n705_));
  AND      g0689(.a(new_n705_), .b(i_2_3_143_0), .O(new_n706_));
  OR       g0690(.a(new_n706_), .b(new_n697_), .O(new_n707_));
  AND      g0691(.a(new_n707_), .b(i_2_3_68_0), .O(new_n708_));
  OR       g0692(.a(i_2_3_86_0), .b(i_2_3_72_0), .O(new_n709_));
  OR       g0693(.a(new_n709_), .b(new_n212_), .O(new_n710_));
  AND      g0694(.a(new_n710_), .b(new_n469_), .O(new_n711_));
  AND      g0695(.a(new_n355_), .b(new_n147_), .O(new_n712_));
  OR       g0696(.a(new_n712_), .b(new_n711_), .O(new_n713_));
  AND      g0697(.a(new_n713_), .b(new_n19_), .O(new_n714_));
  AND      g0698(.a(i_2_3_143_0), .b(i_2_3_79_0), .O(new_n715_));
  AND      g0699(.a(new_n715_), .b(i_2_3_68_0), .O(new_n716_));
  OR       g0700(.a(new_n716_), .b(new_n178_), .O(new_n717_));
  AND      g0701(.a(new_n717_), .b(new_n374_), .O(new_n718_));
  OR       g0702(.a(new_n718_), .b(new_n714_), .O(new_n719_));
  AND      g0703(.a(new_n719_), .b(i_2_3_55_0), .O(new_n720_));
  AND      g0704(.a(new_n374_), .b(i_2_3_79_0), .O(new_n721_));
  AND      g0705(.a(new_n721_), .b(new_n223_), .O(new_n722_));
  OR       g0706(.a(new_n564_), .b(i_2_3_86_0), .O(new_n723_));
  OR       g0707(.a(new_n723_), .b(new_n722_), .O(new_n724_));
  AND      g0708(.a(new_n724_), .b(new_n19_), .O(new_n725_));
  OR       g0709(.a(new_n18_), .b(i_2_3_79_0), .O(new_n726_));
  NAND     g0710(.a(new_n483_), .b(i_2_3_86_0), .O(new_n727_));
  NAND     g0711(.a(new_n727_), .b(new_n726_), .O(new_n728_));
  AND      g0712(.a(new_n728_), .b(new_n77_), .O(new_n729_));
  NAND     g0713(.a(new_n439_), .b(new_n414_), .O(new_n730_));
  OR       g0714(.a(new_n730_), .b(new_n729_), .O(new_n731_));
  OR       g0715(.a(new_n731_), .b(new_n725_), .O(new_n732_));
  AND      g0716(.a(new_n732_), .b(new_n31_), .O(new_n733_));
  OR       g0717(.a(new_n733_), .b(new_n720_), .O(new_n734_));
  OR       g0718(.a(new_n734_), .b(new_n708_), .O(new_n735_));
  AND      g0719(.a(new_n735_), .b(i_2_3_91_0), .O(new_n736_));
  OR       g0720(.a(new_n736_), .b(new_n696_), .O(new_n737_));
  AND      g0721(.a(new_n737_), .b(new_n20_), .O(new_n738_));
  AND      g0722(.a(new_n40_), .b(i_2_3_55_0), .O(new_n739_));
  OR       g0723(.a(new_n739_), .b(new_n353_), .O(new_n740_));
  AND      g0724(.a(new_n740_), .b(new_n77_), .O(new_n741_));
  OR       g0725(.a(new_n40_), .b(i_2_3_68_0), .O(new_n742_));
  AND      g0726(.a(new_n223_), .b(i_2_3_55_0), .O(new_n743_));
  OR       g0727(.a(new_n743_), .b(new_n353_), .O(new_n744_));
  AND      g0728(.a(new_n744_), .b(new_n742_), .O(new_n745_));
  OR       g0729(.a(new_n745_), .b(new_n741_), .O(new_n746_));
  AND      g0730(.a(new_n746_), .b(i_2_3_86_0), .O(new_n747_));
  AND      g0731(.a(new_n458_), .b(new_n213_), .O(new_n748_));
  OR       g0732(.a(new_n748_), .b(new_n747_), .O(new_n749_));
  AND      g0733(.a(new_n749_), .b(i_2_3_91_0), .O(new_n750_));
  AND      g0734(.a(new_n743_), .b(new_n179_), .O(new_n751_));
  OR       g0735(.a(new_n751_), .b(new_n750_), .O(new_n752_));
  AND      g0736(.a(new_n752_), .b(i_2_3_72_0), .O(new_n753_));
  OR       g0737(.a(new_n753_), .b(new_n163_), .O(new_n754_));
  AND      g0738(.a(new_n754_), .b(new_n633_), .O(new_n755_));
  AND      g0739(.a(new_n468_), .b(i_2_3_55_0), .O(new_n756_));
  AND      g0740(.a(new_n756_), .b(new_n625_), .O(new_n757_));
  AND      g0741(.a(new_n757_), .b(new_n163_), .O(new_n758_));
  OR       g0742(.a(new_n758_), .b(new_n755_), .O(new_n759_));
  OR       g0743(.a(new_n759_), .b(new_n738_), .O(new_n760_));
  OR       g0744(.a(new_n760_), .b(new_n682_), .O(new_n761_));
  AND      g0745(.a(new_n761_), .b(i_2_3_29_0), .O(new_n762_));
  AND      g0746(.a(new_n468_), .b(new_n63_), .O(new_n763_));
  OR       g0747(.a(new_n763_), .b(new_n19_), .O(new_n764_));
  OR       g0748(.a(new_n374_), .b(new_n21_), .O(new_n765_));
  AND      g0749(.a(new_n765_), .b(new_n53_), .O(new_n766_));
  OR       g0750(.a(new_n483_), .b(new_n348_), .O(new_n767_));
  AND      g0751(.a(new_n767_), .b(new_n77_), .O(new_n768_));
  OR       g0752(.a(new_n768_), .b(new_n766_), .O(new_n769_));
  OR       g0753(.a(new_n769_), .b(new_n764_), .O(new_n770_));
  AND      g0754(.a(new_n770_), .b(i_2_3_86_0), .O(new_n771_));
  AND      g0755(.a(new_n369_), .b(i_2_3_99_0), .O(new_n772_));
  AND      g0756(.a(new_n511_), .b(i_2_3_72_0), .O(new_n773_));
  OR       g0757(.a(new_n533_), .b(new_n773_), .O(new_n774_));
  OR       g0758(.a(new_n774_), .b(new_n772_), .O(new_n775_));
  AND      g0759(.a(new_n775_), .b(new_n53_), .O(new_n776_));
  OR       g0760(.a(new_n18_), .b(i_2_3_99_0), .O(new_n777_));
  OR       g0761(.a(new_n777_), .b(new_n25_), .O(new_n778_));
  OR       g0762(.a(new_n778_), .b(new_n627_), .O(new_n779_));
  OR       g0763(.a(i_2_3_77_0), .b(i_2_3_68_0), .O(new_n780_));
  OR       g0764(.a(new_n223_), .b(i_2_3_42_0), .O(new_n781_));
  AND      g0765(.a(new_n781_), .b(new_n780_), .O(new_n782_));
  AND      g0766(.a(new_n510_), .b(i_2_3_43_0), .O(new_n783_));
  NAND     g0767(.a(new_n783_), .b(new_n642_), .O(new_n784_));
  OR       g0768(.a(new_n784_), .b(new_n782_), .O(new_n785_));
  NAND     g0769(.a(new_n785_), .b(new_n779_), .O(new_n786_));
  OR       g0770(.a(new_n786_), .b(new_n776_), .O(new_n787_));
  OR       g0771(.a(new_n787_), .b(new_n771_), .O(new_n788_));
  AND      g0772(.a(new_n788_), .b(i_2_3_55_0), .O(new_n789_));
  OR       g0773(.a(new_n539_), .b(new_n348_), .O(new_n790_));
  AND      g0774(.a(new_n790_), .b(new_n194_), .O(new_n791_));
  OR       g0775(.a(new_n468_), .b(i_2_3_72_0), .O(new_n792_));
  NAND     g0776(.a(i_2_3_72_0), .b(i_2_3_68_0), .O(new_n793_));
  NAND     g0777(.a(new_n793_), .b(i_2_3_77_0), .O(new_n794_));
  AND      g0778(.a(new_n794_), .b(new_n236_), .O(new_n795_));
  AND      g0779(.a(new_n795_), .b(new_n792_), .O(new_n796_));
  OR       g0780(.a(new_n796_), .b(new_n791_), .O(new_n797_));
  AND      g0781(.a(new_n797_), .b(i_2_3_86_0), .O(new_n798_));
  OR       g0782(.a(i_2_3_72_0), .b(i_2_3_42_0), .O(new_n799_));
  NOT      g0783(.a(new_n799_), .O(new_n800_));
  OR       g0784(.a(new_n800_), .b(new_n539_), .O(new_n801_));
  AND      g0785(.a(new_n801_), .b(new_n647_), .O(new_n802_));
  OR       g0786(.a(new_n802_), .b(new_n798_), .O(new_n803_));
  OR       g0787(.a(new_n803_), .b(new_n789_), .O(new_n804_));
  AND      g0788(.a(new_n804_), .b(i_2_3_91_0), .O(new_n805_));
  AND      g0789(.a(new_n533_), .b(new_n128_), .O(new_n806_));
  AND      g0790(.a(new_n212_), .b(new_n22_), .O(new_n807_));
  AND      g0791(.a(new_n807_), .b(new_n806_), .O(new_n808_));
  NAND     g0792(.a(new_n192_), .b(i_2_3_77_0), .O(new_n809_));
  AND      g0793(.a(new_n809_), .b(new_n53_), .O(new_n810_));
  AND      g0794(.a(new_n715_), .b(new_n381_), .O(new_n811_));
  OR       g0795(.a(new_n811_), .b(new_n810_), .O(new_n812_));
  AND      g0796(.a(new_n812_), .b(i_2_3_72_0), .O(new_n813_));
  AND      g0797(.a(new_n525_), .b(new_n25_), .O(new_n814_));
  AND      g0798(.a(new_n549_), .b(new_n70_), .O(new_n815_));
  OR       g0799(.a(new_n815_), .b(new_n814_), .O(new_n816_));
  OR       g0800(.a(new_n816_), .b(new_n813_), .O(new_n817_));
  AND      g0801(.a(new_n817_), .b(i_2_3_68_0), .O(new_n818_));
  NAND     g0802(.a(new_n237_), .b(new_n40_), .O(new_n819_));
  OR       g0803(.a(i_2_3_72_0), .b(new_n53_), .O(new_n820_));
  AND      g0804(.a(new_n820_), .b(new_n633_), .O(new_n821_));
  AND      g0805(.a(new_n821_), .b(new_n819_), .O(new_n822_));
  OR       g0806(.a(new_n822_), .b(new_n818_), .O(new_n823_));
  AND      g0807(.a(new_n823_), .b(new_n56_), .O(new_n824_));
  OR       g0808(.a(new_n824_), .b(new_n808_), .O(new_n825_));
  OR       g0809(.a(new_n825_), .b(new_n805_), .O(new_n826_));
  AND      g0810(.a(new_n826_), .b(new_n20_), .O(new_n827_));
  AND      g0811(.a(new_n533_), .b(new_n53_), .O(new_n828_));
  AND      g0812(.a(new_n399_), .b(new_n395_), .O(new_n829_));
  OR       g0813(.a(new_n829_), .b(new_n84_), .O(new_n830_));
  AND      g0814(.a(new_n830_), .b(new_n828_), .O(new_n831_));
  NOT      g0815(.a(new_n701_), .O(new_n832_));
  NOT      g0816(.a(new_n782_), .O(new_n833_));
  AND      g0817(.a(new_n833_), .b(new_n30_), .O(new_n834_));
  AND      g0818(.a(new_n834_), .b(new_n832_), .O(new_n835_));
  OR       g0819(.a(new_n835_), .b(new_n831_), .O(new_n836_));
  AND      g0820(.a(new_n836_), .b(i_2_3_91_0), .O(new_n837_));
  OR       g0821(.a(new_n837_), .b(new_n827_), .O(new_n838_));
  AND      g0822(.a(new_n838_), .b(new_n31_), .O(new_n839_));
  AND      g0823(.a(new_n533_), .b(new_n77_), .O(new_n840_));
  AND      g0824(.a(new_n430_), .b(new_n99_), .O(new_n841_));
  OR       g0825(.a(new_n841_), .b(new_n575_), .O(new_n842_));
  AND      g0826(.a(new_n842_), .b(new_n53_), .O(new_n843_));
  OR       g0827(.a(new_n843_), .b(new_n840_), .O(new_n844_));
  AND      g0828(.a(new_n844_), .b(new_n21_), .O(new_n845_));
  OR       g0829(.a(i_2_3_143_0), .b(new_n25_), .O(new_n846_));
  AND      g0830(.a(i_2_3_79_0), .b(i_2_3_68_0), .O(new_n847_));
  AND      g0831(.a(new_n847_), .b(new_n846_), .O(new_n848_));
  OR       g0832(.a(new_n19_), .b(i_2_3_72_0), .O(new_n849_));
  AND      g0833(.a(new_n849_), .b(new_n341_), .O(new_n850_));
  AND      g0834(.a(new_n850_), .b(new_n848_), .O(new_n851_));
  OR       g0835(.a(new_n851_), .b(new_n845_), .O(new_n852_));
  AND      g0836(.a(new_n852_), .b(new_n20_), .O(new_n853_));
  AND      g0837(.a(new_n533_), .b(new_n352_), .O(new_n854_));
  OR       g0838(.a(new_n854_), .b(new_n853_), .O(new_n855_));
  AND      g0839(.a(new_n855_), .b(i_2_3_99_0), .O(new_n856_));
  NOT      g0840(.a(new_n94_), .O(new_n857_));
  NOT      g0841(.a(new_n793_), .O(new_n858_));
  AND      g0842(.a(new_n858_), .b(new_n857_), .O(new_n859_));
  AND      g0843(.a(new_n859_), .b(new_n326_), .O(new_n860_));
  OR       g0844(.a(new_n860_), .b(new_n856_), .O(new_n861_));
  AND      g0845(.a(new_n861_), .b(i_2_3_91_0), .O(new_n862_));
  AND      g0846(.a(new_n854_), .b(new_n305_), .O(new_n863_));
  OR       g0847(.a(new_n863_), .b(new_n862_), .O(new_n864_));
  AND      g0848(.a(new_n864_), .b(i_2_3_55_0), .O(new_n865_));
  AND      g0849(.a(new_n715_), .b(new_n154_), .O(new_n866_));
  AND      g0850(.a(new_n866_), .b(new_n41_), .O(new_n867_));
  AND      g0851(.a(new_n867_), .b(new_n806_), .O(new_n868_));
  OR       g0852(.a(new_n868_), .b(new_n865_), .O(new_n869_));
  OR       g0853(.a(new_n869_), .b(new_n839_), .O(new_n870_));
  OR       g0854(.a(new_n870_), .b(new_n762_), .O(new_n871_));
  OR       g0855(.a(new_n871_), .b(new_n524_), .O(new_n872_));
  AND      g0856(.a(new_n872_), .b(new_n17_), .O(new_n873_));
  AND      g0857(.a(new_n18_), .b(i_2_3_79_0), .O(new_n874_));
  OR       g0858(.a(new_n17_), .b(i_2_3_29_0), .O(new_n875_));
  OR       g0859(.a(new_n875_), .b(i_2_3_55_0), .O(new_n876_));
  NAND     g0860(.a(new_n876_), .b(new_n40_), .O(new_n877_));
  AND      g0861(.a(new_n877_), .b(new_n874_), .O(new_n878_));
  AND      g0862(.a(new_n777_), .b(i_2_3_29_0), .O(new_n879_));
  AND      g0863(.a(new_n879_), .b(new_n21_), .O(new_n880_));
  OR       g0864(.a(new_n880_), .b(new_n20_), .O(new_n881_));
  AND      g0865(.a(new_n881_), .b(new_n206_), .O(new_n882_));
  OR       g0866(.a(new_n882_), .b(new_n878_), .O(new_n883_));
  AND      g0867(.a(new_n883_), .b(i_2_3_72_0), .O(new_n884_));
  NAND     g0868(.a(new_n875_), .b(i_2_3_79_0), .O(new_n885_));
  AND      g0869(.a(i_2_3_99_0), .b(new_n25_), .O(new_n886_));
  AND      g0870(.a(new_n886_), .b(new_n885_), .O(new_n887_));
  OR       g0871(.a(new_n887_), .b(new_n857_), .O(new_n888_));
  AND      g0872(.a(new_n888_), .b(new_n18_), .O(new_n889_));
  OR       g0873(.a(new_n889_), .b(new_n884_), .O(new_n890_));
  AND      g0874(.a(new_n890_), .b(new_n19_), .O(new_n891_));
  AND      g0875(.a(i_2_3_72_0), .b(i_2_3_29_0), .O(new_n892_));
  AND      g0876(.a(new_n374_), .b(new_n18_), .O(new_n893_));
  OR       g0877(.a(new_n893_), .b(new_n892_), .O(new_n894_));
  NAND     g0878(.a(new_n846_), .b(new_n40_), .O(new_n895_));
  AND      g0879(.a(new_n895_), .b(new_n21_), .O(new_n896_));
  OR       g0880(.a(new_n896_), .b(new_n894_), .O(new_n897_));
  AND      g0881(.a(new_n897_), .b(new_n267_), .O(new_n898_));
  OR       g0882(.a(new_n898_), .b(new_n891_), .O(new_n899_));
  AND      g0883(.a(new_n899_), .b(i_2_3_86_0), .O(new_n900_));
  AND      g0884(.a(new_n18_), .b(i_2_3_29_0), .O(new_n901_));
  OR       g0885(.a(new_n901_), .b(new_n212_), .O(new_n902_));
  AND      g0886(.a(new_n902_), .b(new_n369_), .O(new_n903_));
  OR       g0887(.a(i_2_3_143_0), .b(i_2_3_72_0), .O(new_n904_));
  NAND     g0888(.a(new_n904_), .b(i_2_3_79_0), .O(new_n905_));
  AND      g0889(.a(new_n905_), .b(i_2_3_77_0), .O(new_n906_));
  OR       g0890(.a(i_2_3_143_0), .b(i_2_3_79_0), .O(new_n907_));
  AND      g0891(.a(new_n18_), .b(i_2_3_43_0), .O(new_n908_));
  NOT      g0892(.a(new_n908_), .O(new_n909_));
  AND      g0893(.a(new_n909_), .b(new_n40_), .O(new_n910_));
  NAND     g0894(.a(new_n910_), .b(new_n907_), .O(new_n911_));
  OR       g0895(.a(new_n911_), .b(new_n906_), .O(new_n912_));
  AND      g0896(.a(new_n912_), .b(i_2_3_29_0), .O(new_n913_));
  OR       g0897(.a(new_n913_), .b(new_n903_), .O(new_n914_));
  AND      g0898(.a(new_n914_), .b(new_n20_), .O(new_n915_));
  OR       g0899(.a(new_n915_), .b(new_n900_), .O(new_n916_));
  AND      g0900(.a(new_n916_), .b(i_2_3_68_0), .O(new_n917_));
  OR       g0901(.a(new_n632_), .b(i_2_3_143_0), .O(new_n918_));
  NOT      g0902(.a(new_n918_), .O(new_n919_));
  AND      g0903(.a(new_n919_), .b(new_n305_), .O(new_n920_));
  AND      g0904(.a(new_n920_), .b(i_2_3_86_0), .O(new_n921_));
  OR       g0905(.a(new_n355_), .b(new_n193_), .O(new_n922_));
  AND      g0906(.a(new_n922_), .b(i_2_3_72_0), .O(new_n923_));
  NAND     g0907(.a(new_n303_), .b(i_2_3_79_0), .O(new_n924_));
  AND      g0908(.a(new_n924_), .b(new_n400_), .O(new_n925_));
  OR       g0909(.a(new_n925_), .b(new_n923_), .O(new_n926_));
  AND      g0910(.a(new_n926_), .b(new_n19_), .O(new_n927_));
  AND      g0911(.a(i_2_3_142_0), .b(i_2_3_77_0), .O(new_n928_));
  OR       g0912(.a(new_n928_), .b(i_2_3_72_0), .O(new_n929_));
  AND      g0913(.a(new_n929_), .b(new_n381_), .O(new_n930_));
  AND      g0914(.a(new_n626_), .b(new_n21_), .O(new_n931_));
  OR       g0915(.a(new_n931_), .b(new_n575_), .O(new_n932_));
  OR       g0916(.a(new_n932_), .b(new_n930_), .O(new_n933_));
  AND      g0917(.a(new_n933_), .b(new_n18_), .O(new_n934_));
  OR       g0918(.a(new_n934_), .b(new_n927_), .O(new_n935_));
  AND      g0919(.a(new_n935_), .b(new_n20_), .O(new_n936_));
  AND      g0920(.a(new_n212_), .b(new_n18_), .O(new_n937_));
  AND      g0921(.a(new_n340_), .b(i_2_3_77_0), .O(new_n938_));
  AND      g0922(.a(new_n938_), .b(new_n937_), .O(new_n939_));
  OR       g0923(.a(new_n939_), .b(new_n936_), .O(new_n940_));
  AND      g0924(.a(new_n940_), .b(i_2_3_29_0), .O(new_n941_));
  OR       g0925(.a(new_n941_), .b(new_n921_), .O(new_n942_));
  OR       g0926(.a(new_n942_), .b(new_n917_), .O(new_n943_));
  AND      g0927(.a(new_n943_), .b(new_n53_), .O(new_n944_));
  AND      g0928(.a(new_n575_), .b(new_n40_), .O(new_n945_));
  OR       g0929(.a(new_n19_), .b(i_2_3_43_0), .O(new_n946_));
  AND      g0930(.a(new_n946_), .b(i_2_3_29_0), .O(new_n947_));
  AND      g0931(.a(new_n20_), .b(i_2_3_68_0), .O(new_n948_));
  OR       g0932(.a(new_n948_), .b(new_n947_), .O(new_n949_));
  OR       g0933(.a(new_n949_), .b(new_n945_), .O(new_n950_));
  AND      g0934(.a(new_n950_), .b(new_n21_), .O(new_n951_));
  AND      g0935(.a(i_2_3_142_0), .b(new_n223_), .O(new_n952_));
  AND      g0936(.a(new_n952_), .b(new_n525_), .O(new_n953_));
  AND      g0937(.a(new_n105_), .b(new_n40_), .O(new_n954_));
  OR       g0938(.a(new_n954_), .b(new_n953_), .O(new_n955_));
  AND      g0939(.a(new_n955_), .b(new_n77_), .O(new_n956_));
  AND      g0940(.a(i_2_3_68_0), .b(i_2_3_29_0), .O(new_n957_));
  AND      g0941(.a(new_n957_), .b(new_n525_), .O(new_n958_));
  OR       g0942(.a(new_n633_), .b(new_n533_), .O(new_n959_));
  OR       g0943(.a(new_n959_), .b(new_n378_), .O(new_n960_));
  AND      g0944(.a(new_n960_), .b(new_n20_), .O(new_n961_));
  OR       g0945(.a(new_n961_), .b(new_n958_), .O(new_n962_));
  OR       g0946(.a(new_n962_), .b(new_n956_), .O(new_n963_));
  OR       g0947(.a(new_n963_), .b(new_n951_), .O(new_n964_));
  AND      g0948(.a(new_n964_), .b(i_2_3_72_0), .O(new_n965_));
  AND      g0949(.a(new_n40_), .b(i_2_3_43_0), .O(new_n966_));
  OR       g0950(.a(new_n966_), .b(new_n20_), .O(new_n967_));
  AND      g0951(.a(new_n967_), .b(i_2_3_29_0), .O(new_n968_));
  OR       g0952(.a(new_n647_), .b(new_n301_), .O(new_n969_));
  AND      g0953(.a(new_n969_), .b(new_n25_), .O(new_n970_));
  OR       g0954(.a(new_n970_), .b(new_n968_), .O(new_n971_));
  AND      g0955(.a(new_n971_), .b(new_n19_), .O(new_n972_));
  AND      g0956(.a(new_n742_), .b(i_2_3_29_0), .O(new_n973_));
  OR       g0957(.a(new_n952_), .b(i_2_3_99_0), .O(new_n974_));
  AND      g0958(.a(new_n974_), .b(new_n973_), .O(new_n975_));
  OR       g0959(.a(new_n948_), .b(new_n647_), .O(new_n976_));
  OR       g0960(.a(new_n976_), .b(new_n975_), .O(new_n977_));
  AND      g0961(.a(new_n977_), .b(i_2_3_86_0), .O(new_n978_));
  OR       g0962(.a(new_n978_), .b(new_n972_), .O(new_n979_));
  OR       g0963(.a(new_n979_), .b(new_n965_), .O(new_n980_));
  AND      g0964(.a(new_n980_), .b(new_n18_), .O(new_n981_));
  NAND     g0965(.a(new_n892_), .b(i_2_3_99_0), .O(new_n982_));
  OR       g0966(.a(new_n875_), .b(new_n709_), .O(new_n983_));
  NAND     g0967(.a(new_n983_), .b(new_n982_), .O(new_n984_));
  AND      g0968(.a(new_n984_), .b(i_2_3_68_0), .O(new_n985_));
  AND      g0969(.a(new_n303_), .b(new_n267_), .O(new_n986_));
  AND      g0970(.a(new_n105_), .b(new_n44_), .O(new_n987_));
  OR       g0971(.a(new_n987_), .b(new_n986_), .O(new_n988_));
  OR       g0972(.a(new_n988_), .b(new_n985_), .O(new_n989_));
  AND      g0973(.a(new_n989_), .b(new_n19_), .O(new_n990_));
  AND      g0974(.a(new_n301_), .b(i_2_3_68_0), .O(new_n991_));
  OR       g0975(.a(new_n374_), .b(i_2_3_68_0), .O(new_n992_));
  AND      g0976(.a(new_n992_), .b(new_n20_), .O(new_n993_));
  AND      g0977(.a(new_n973_), .b(new_n431_), .O(new_n994_));
  OR       g0978(.a(new_n994_), .b(new_n993_), .O(new_n995_));
  AND      g0979(.a(new_n995_), .b(i_2_3_86_0), .O(new_n996_));
  OR       g0980(.a(new_n996_), .b(new_n991_), .O(new_n997_));
  OR       g0981(.a(new_n997_), .b(new_n990_), .O(new_n998_));
  AND      g0982(.a(new_n998_), .b(new_n21_), .O(new_n999_));
  OR       g0983(.a(new_n533_), .b(new_n381_), .O(new_n1000_));
  AND      g0984(.a(new_n1000_), .b(new_n794_), .O(new_n1001_));
  OR       g0985(.a(new_n305_), .b(new_n196_), .O(new_n1002_));
  OR       g0986(.a(new_n1002_), .b(new_n1001_), .O(new_n1003_));
  AND      g0987(.a(new_n1003_), .b(i_2_3_86_0), .O(new_n1004_));
  AND      g0988(.a(new_n948_), .b(new_n77_), .O(new_n1005_));
  OR       g0989(.a(new_n1005_), .b(new_n1004_), .O(new_n1006_));
  AND      g0990(.a(new_n1006_), .b(i_2_3_29_0), .O(new_n1007_));
  OR       g0991(.a(new_n458_), .b(new_n178_), .O(new_n1008_));
  AND      g0992(.a(new_n1008_), .b(new_n19_), .O(new_n1009_));
  OR       g0993(.a(new_n1009_), .b(new_n459_), .O(new_n1010_));
  AND      g0994(.a(new_n1010_), .b(new_n20_), .O(new_n1011_));
  OR       g0995(.a(new_n1011_), .b(new_n1007_), .O(new_n1012_));
  OR       g0996(.a(new_n1012_), .b(new_n999_), .O(new_n1013_));
  OR       g0997(.a(new_n1013_), .b(new_n981_), .O(new_n1014_));
  AND      g0998(.a(new_n1014_), .b(new_n53_), .O(new_n1015_));
  OR       g0999(.a(i_2_3_138_0), .b(i_2_3_77_0), .O(new_n1016_));
  OR       g1000(.a(new_n709_), .b(new_n17_), .O(new_n1017_));
  NAND     g1001(.a(new_n1017_), .b(new_n1016_), .O(new_n1018_));
  AND      g1002(.a(new_n18_), .b(i_2_3_99_0), .O(new_n1019_));
  AND      g1003(.a(new_n1019_), .b(new_n511_), .O(new_n1020_));
  AND      g1004(.a(new_n1020_), .b(new_n1018_), .O(new_n1021_));
  OR       g1005(.a(new_n918_), .b(new_n481_), .O(new_n1022_));
  OR       g1006(.a(i_2_3_143_0), .b(i_2_3_77_0), .O(new_n1023_));
  NOT      g1007(.a(new_n1023_), .O(new_n1024_));
  AND      g1008(.a(new_n546_), .b(new_n21_), .O(new_n1025_));
  OR       g1009(.a(new_n1025_), .b(new_n1019_), .O(new_n1026_));
  OR       g1010(.a(new_n1026_), .b(new_n1024_), .O(new_n1027_));
  AND      g1011(.a(new_n1027_), .b(i_2_3_72_0), .O(new_n1028_));
  OR       g1012(.a(new_n1028_), .b(new_n625_), .O(new_n1029_));
  AND      g1013(.a(new_n1029_), .b(i_2_3_68_0), .O(new_n1030_));
  AND      g1014(.a(new_n549_), .b(i_2_3_68_0), .O(new_n1031_));
  AND      g1015(.a(new_n1031_), .b(new_n1026_), .O(new_n1032_));
  NAND     g1016(.a(new_n1023_), .b(new_n311_), .O(new_n1033_));
  AND      g1017(.a(new_n546_), .b(i_2_3_99_0), .O(new_n1034_));
  AND      g1018(.a(new_n1034_), .b(new_n1033_), .O(new_n1035_));
  OR       g1019(.a(new_n1035_), .b(new_n1032_), .O(new_n1036_));
  OR       g1020(.a(new_n1036_), .b(new_n1030_), .O(new_n1037_));
  NAND     g1021(.a(new_n1037_), .b(new_n20_), .O(new_n1038_));
  NAND     g1022(.a(new_n1038_), .b(new_n1022_), .O(new_n1039_));
  AND      g1023(.a(new_n1039_), .b(i_2_3_86_0), .O(new_n1040_));
  OR       g1024(.a(new_n1040_), .b(new_n1021_), .O(new_n1041_));
  OR       g1025(.a(new_n1041_), .b(new_n1015_), .O(new_n1042_));
  AND      g1026(.a(new_n1042_), .b(i_2_3_55_0), .O(new_n1043_));
  AND      g1027(.a(new_n921_), .b(i_2_3_68_0), .O(new_n1044_));
  AND      g1028(.a(new_n1024_), .b(new_n765_), .O(new_n1045_));
  OR       g1029(.a(new_n1045_), .b(new_n1030_), .O(new_n1046_));
  AND      g1030(.a(new_n1046_), .b(new_n20_), .O(new_n1047_));
  NOT      g1031(.a(new_n780_), .O(new_n1048_));
  AND      g1032(.a(new_n937_), .b(new_n1048_), .O(new_n1049_));
  OR       g1033(.a(new_n1049_), .b(new_n565_), .O(new_n1050_));
  AND      g1034(.a(new_n1050_), .b(new_n77_), .O(new_n1051_));
  OR       g1035(.a(new_n1051_), .b(new_n1047_), .O(new_n1052_));
  AND      g1036(.a(new_n1052_), .b(i_2_3_86_0), .O(new_n1053_));
  NOT      g1037(.a(new_n715_), .O(new_n1054_));
  NAND     g1038(.a(new_n907_), .b(i_2_3_138_0), .O(new_n1055_));
  AND      g1039(.a(new_n1055_), .b(new_n1054_), .O(new_n1056_));
  OR       g1040(.a(new_n948_), .b(new_n305_), .O(new_n1057_));
  OR       g1041(.a(new_n1057_), .b(new_n893_), .O(new_n1058_));
  OR       g1042(.a(new_n1058_), .b(new_n462_), .O(new_n1059_));
  OR       g1043(.a(new_n1059_), .b(new_n1056_), .O(new_n1060_));
  AND      g1044(.a(new_n1060_), .b(new_n19_), .O(new_n1061_));
  AND      g1045(.a(new_n948_), .b(new_n778_), .O(new_n1062_));
  OR       g1046(.a(new_n1062_), .b(new_n21_), .O(new_n1063_));
  OR       g1047(.a(i_2_3_143_0), .b(i_2_3_68_0), .O(new_n1064_));
  NOT      g1048(.a(new_n1064_), .O(new_n1065_));
  OR       g1049(.a(new_n1065_), .b(new_n1019_), .O(new_n1066_));
  OR       g1050(.a(new_n1066_), .b(new_n993_), .O(new_n1067_));
  AND      g1051(.a(new_n1067_), .b(new_n1063_), .O(new_n1068_));
  OR       g1052(.a(new_n1068_), .b(new_n1061_), .O(new_n1069_));
  AND      g1053(.a(new_n1069_), .b(i_2_3_86_0), .O(new_n1070_));
  AND      g1054(.a(new_n721_), .b(i_2_3_43_0), .O(new_n1071_));
  OR       g1055(.a(new_n1071_), .b(new_n513_), .O(new_n1072_));
  AND      g1056(.a(new_n1072_), .b(new_n18_), .O(new_n1073_));
  OR       g1057(.a(new_n1073_), .b(new_n647_), .O(new_n1074_));
  AND      g1058(.a(new_n1074_), .b(new_n20_), .O(new_n1075_));
  AND      g1059(.a(new_n642_), .b(new_n20_), .O(new_n1076_));
  OR       g1060(.a(i_2_3_79_0), .b(new_n223_), .O(new_n1077_));
  NAND     g1061(.a(new_n846_), .b(new_n1077_), .O(new_n1078_));
  AND      g1062(.a(new_n1078_), .b(new_n1076_), .O(new_n1079_));
  AND      g1063(.a(new_n1076_), .b(new_n147_), .O(new_n1080_));
  OR       g1064(.a(new_n1080_), .b(new_n77_), .O(new_n1081_));
  AND      g1065(.a(new_n1055_), .b(i_2_3_99_0), .O(new_n1082_));
  AND      g1066(.a(new_n1082_), .b(new_n1081_), .O(new_n1083_));
  OR       g1067(.a(new_n1083_), .b(new_n1079_), .O(new_n1084_));
  AND      g1068(.a(new_n1084_), .b(new_n19_), .O(new_n1085_));
  OR       g1069(.a(new_n1085_), .b(new_n1075_), .O(new_n1086_));
  OR       g1070(.a(new_n1086_), .b(new_n1070_), .O(new_n1087_));
  AND      g1071(.a(new_n1087_), .b(i_2_3_55_0), .O(new_n1088_));
  OR       g1072(.a(new_n1088_), .b(new_n920_), .O(new_n1089_));
  OR       g1073(.a(new_n1089_), .b(new_n1053_), .O(new_n1090_));
  AND      g1074(.a(new_n1090_), .b(i_2_3_29_0), .O(new_n1091_));
  OR       g1075(.a(new_n1091_), .b(new_n1044_), .O(new_n1092_));
  OR       g1076(.a(new_n1092_), .b(new_n1043_), .O(new_n1093_));
  OR       g1077(.a(new_n1093_), .b(new_n944_), .O(new_n1094_));
  AND      g1078(.a(new_n1094_), .b(new_n31_), .O(new_n1095_));
  NOT      g1079(.a(new_n726_), .O(new_n1096_));
  AND      g1080(.a(new_n892_), .b(new_n1096_), .O(new_n1097_));
  OR       g1081(.a(new_n1019_), .b(new_n147_), .O(new_n1098_));
  AND      g1082(.a(new_n1098_), .b(new_n879_), .O(new_n1099_));
  OR       g1083(.a(new_n1099_), .b(new_n253_), .O(new_n1100_));
  AND      g1084(.a(new_n1100_), .b(new_n957_), .O(new_n1101_));
  AND      g1085(.a(new_n715_), .b(i_2_3_142_0), .O(new_n1102_));
  OR       g1086(.a(new_n1102_), .b(new_n511_), .O(new_n1103_));
  AND      g1087(.a(new_n1103_), .b(i_2_3_72_0), .O(new_n1104_));
  AND      g1088(.a(new_n21_), .b(i_2_3_29_0), .O(new_n1105_));
  AND      g1089(.a(new_n1105_), .b(new_n909_), .O(new_n1106_));
  OR       g1090(.a(new_n1106_), .b(new_n1104_), .O(new_n1107_));
  AND      g1091(.a(new_n1107_), .b(i_2_3_99_0), .O(new_n1108_));
  OR       g1092(.a(new_n1108_), .b(new_n1101_), .O(new_n1109_));
  AND      g1093(.a(new_n1109_), .b(new_n19_), .O(new_n1110_));
  OR       g1094(.a(new_n1110_), .b(new_n1097_), .O(new_n1111_));
  AND      g1095(.a(new_n1111_), .b(new_n53_), .O(new_n1112_));
  OR       g1096(.a(new_n381_), .b(new_n18_), .O(new_n1113_));
  AND      g1097(.a(new_n1113_), .b(i_2_3_29_0), .O(new_n1114_));
  AND      g1098(.a(new_n905_), .b(i_2_3_99_0), .O(new_n1115_));
  OR       g1099(.a(new_n1115_), .b(new_n1114_), .O(new_n1116_));
  AND      g1100(.a(new_n1116_), .b(i_2_3_68_0), .O(new_n1117_));
  NOT      g1101(.a(new_n459_), .O(new_n1118_));
  OR       g1102(.a(i_2_3_143_0), .b(new_n17_), .O(new_n1119_));
  OR       g1103(.a(new_n1119_), .b(new_n19_), .O(new_n1120_));
  OR       g1104(.a(new_n1120_), .b(new_n278_), .O(new_n1121_));
  NAND     g1105(.a(new_n1121_), .b(new_n1118_), .O(new_n1122_));
  AND      g1106(.a(new_n1122_), .b(i_2_3_43_0), .O(new_n1123_));
  AND      g1107(.a(new_n901_), .b(i_2_3_72_0), .O(new_n1124_));
  OR       g1108(.a(new_n1124_), .b(new_n1123_), .O(new_n1125_));
  OR       g1109(.a(new_n1125_), .b(new_n1117_), .O(new_n1126_));
  AND      g1110(.a(new_n1126_), .b(new_n53_), .O(new_n1127_));
  AND      g1111(.a(new_n901_), .b(new_n467_), .O(new_n1128_));
  AND      g1112(.a(new_n1128_), .b(new_n464_), .O(new_n1129_));
  AND      g1113(.a(new_n894_), .b(new_n21_), .O(new_n1130_));
  OR       g1114(.a(new_n1130_), .b(new_n1099_), .O(new_n1131_));
  AND      g1115(.a(new_n1131_), .b(i_2_3_68_0), .O(new_n1132_));
  AND      g1116(.a(new_n1128_), .b(new_n21_), .O(new_n1133_));
  OR       g1117(.a(new_n1133_), .b(new_n1132_), .O(new_n1134_));
  AND      g1118(.a(new_n1134_), .b(new_n19_), .O(new_n1135_));
  OR       g1119(.a(new_n1135_), .b(new_n1129_), .O(new_n1136_));
  OR       g1120(.a(new_n1136_), .b(new_n1127_), .O(new_n1137_));
  AND      g1121(.a(new_n1137_), .b(i_2_3_86_0), .O(new_n1138_));
  OR       g1122(.a(new_n1138_), .b(new_n1112_), .O(new_n1139_));
  AND      g1123(.a(new_n1139_), .b(i_2_3_55_0), .O(new_n1140_));
  AND      g1124(.a(new_n937_), .b(new_n592_), .O(new_n1141_));
  OR       g1125(.a(new_n1023_), .b(new_n99_), .O(new_n1142_));
  NAND     g1126(.a(new_n1142_), .b(new_n334_), .O(new_n1143_));
  AND      g1127(.a(new_n1143_), .b(new_n77_), .O(new_n1144_));
  AND      g1128(.a(new_n1025_), .b(new_n1023_), .O(new_n1145_));
  OR       g1129(.a(new_n1145_), .b(new_n1144_), .O(new_n1146_));
  AND      g1130(.a(new_n1146_), .b(i_2_3_72_0), .O(new_n1147_));
  AND      g1131(.a(new_n1024_), .b(new_n378_), .O(new_n1148_));
  OR       g1132(.a(new_n1148_), .b(new_n212_), .O(new_n1149_));
  OR       g1133(.a(new_n1149_), .b(new_n1147_), .O(new_n1150_));
  AND      g1134(.a(new_n1150_), .b(i_2_3_68_0), .O(new_n1151_));
  OR       g1135(.a(new_n1151_), .b(new_n1141_), .O(new_n1152_));
  AND      g1136(.a(new_n1152_), .b(new_n53_), .O(new_n1153_));
  AND      g1137(.a(new_n893_), .b(new_n533_), .O(new_n1154_));
  AND      g1138(.a(new_n1154_), .b(new_n139_), .O(new_n1155_));
  OR       g1139(.a(new_n1155_), .b(new_n1153_), .O(new_n1156_));
  AND      g1140(.a(new_n1156_), .b(i_2_3_29_0), .O(new_n1157_));
  NOT      g1141(.a(new_n237_), .O(new_n1158_));
  AND      g1142(.a(new_n874_), .b(new_n1158_), .O(new_n1159_));
  AND      g1143(.a(new_n1159_), .b(new_n828_), .O(new_n1160_));
  OR       g1144(.a(new_n1160_), .b(new_n1157_), .O(new_n1161_));
  OR       g1145(.a(new_n1161_), .b(new_n1140_), .O(new_n1162_));
  AND      g1146(.a(new_n1162_), .b(new_n20_), .O(new_n1163_));
  OR       g1147(.a(new_n20_), .b(i_2_3_72_0), .O(new_n1164_));
  AND      g1148(.a(new_n1164_), .b(new_n18_), .O(new_n1165_));
  OR       g1149(.a(new_n1165_), .b(new_n458_), .O(new_n1166_));
  AND      g1150(.a(new_n1166_), .b(i_2_3_29_0), .O(new_n1167_));
  OR       g1151(.a(new_n1167_), .b(new_n459_), .O(new_n1168_));
  AND      g1152(.a(new_n1168_), .b(new_n21_), .O(new_n1169_));
  AND      g1153(.a(new_n18_), .b(i_2_3_142_0), .O(new_n1170_));
  NAND     g1154(.a(new_n1170_), .b(new_n212_), .O(new_n1171_));
  NOT      g1155(.a(new_n1171_), .O(new_n1172_));
  OR       g1156(.a(new_n1172_), .b(new_n196_), .O(new_n1173_));
  AND      g1157(.a(new_n1173_), .b(new_n359_), .O(new_n1174_));
  OR       g1158(.a(new_n1174_), .b(new_n1020_), .O(new_n1175_));
  AND      g1159(.a(new_n1175_), .b(new_n77_), .O(new_n1176_));
  NOT      g1160(.a(new_n642_), .O(new_n1177_));
  AND      g1161(.a(new_n901_), .b(new_n886_), .O(new_n1178_));
  AND      g1162(.a(new_n1178_), .b(new_n1177_), .O(new_n1179_));
  OR       g1163(.a(new_n1179_), .b(new_n316_), .O(new_n1180_));
  AND      g1164(.a(new_n1180_), .b(i_2_3_142_0), .O(new_n1181_));
  AND      g1165(.a(new_n908_), .b(new_n892_), .O(new_n1182_));
  AND      g1166(.a(new_n948_), .b(new_n147_), .O(new_n1183_));
  OR       g1167(.a(new_n1183_), .b(new_n1182_), .O(new_n1184_));
  OR       g1168(.a(new_n1184_), .b(new_n1181_), .O(new_n1185_));
  OR       g1169(.a(new_n1185_), .b(new_n1176_), .O(new_n1186_));
  OR       g1170(.a(new_n1186_), .b(new_n1169_), .O(new_n1187_));
  AND      g1171(.a(new_n688_), .b(new_n326_), .O(new_n1188_));
  AND      g1172(.a(new_n1188_), .b(new_n1187_), .O(new_n1189_));
  OR       g1173(.a(new_n1189_), .b(new_n1163_), .O(new_n1190_));
  OR       g1174(.a(new_n1190_), .b(new_n1095_), .O(new_n1191_));
  AND      g1175(.a(new_n1191_), .b(i_2_3_91_0), .O(new_n1192_));
  NAND     g1176(.a(new_n1119_), .b(i_2_3_43_0), .O(new_n1193_));
  AND      g1177(.a(new_n1193_), .b(i_2_3_29_0), .O(new_n1194_));
  AND      g1178(.a(i_2_3_142_0), .b(new_n77_), .O(new_n1195_));
  OR       g1179(.a(new_n1195_), .b(i_2_3_55_0), .O(new_n1196_));
  AND      g1180(.a(new_n1196_), .b(i_2_3_68_0), .O(new_n1197_));
  OR       g1181(.a(new_n1197_), .b(new_n1194_), .O(new_n1198_));
  AND      g1182(.a(new_n1198_), .b(i_2_3_72_0), .O(new_n1199_));
  AND      g1183(.a(new_n183_), .b(i_2_3_68_0), .O(new_n1200_));
  OR       g1184(.a(new_n1200_), .b(new_n1199_), .O(new_n1201_));
  AND      g1185(.a(new_n1201_), .b(i_2_3_99_0), .O(new_n1202_));
  AND      g1186(.a(new_n18_), .b(i_2_3_68_0), .O(new_n1203_));
  AND      g1187(.a(new_n1203_), .b(new_n77_), .O(new_n1204_));
  AND      g1188(.a(new_n1204_), .b(new_n183_), .O(new_n1205_));
  OR       g1189(.a(new_n1205_), .b(new_n1202_), .O(new_n1206_));
  AND      g1190(.a(new_n1206_), .b(new_n21_), .O(new_n1207_));
  AND      g1191(.a(new_n957_), .b(new_n893_), .O(new_n1208_));
  OR       g1192(.a(new_n1208_), .b(new_n1207_), .O(new_n1209_));
  AND      g1193(.a(new_n1209_), .b(new_n19_), .O(new_n1210_));
  AND      g1194(.a(new_n886_), .b(new_n874_), .O(new_n1211_));
  AND      g1195(.a(new_n1211_), .b(new_n1200_), .O(new_n1212_));
  OR       g1196(.a(new_n1212_), .b(new_n1210_), .O(new_n1213_));
  AND      g1197(.a(new_n1213_), .b(new_n20_), .O(new_n1214_));
  NOT      g1198(.a(new_n702_), .O(new_n1215_));
  AND      g1199(.a(new_n1172_), .b(new_n1215_), .O(new_n1216_));
  AND      g1200(.a(new_n1216_), .b(new_n1200_), .O(new_n1217_));
  OR       g1201(.a(new_n1217_), .b(new_n1214_), .O(new_n1218_));
  AND      g1202(.a(new_n1218_), .b(i_2_3_86_0), .O(new_n1219_));
  NOT      g1203(.a(new_n627_), .O(new_n1220_));
  NOT      g1204(.a(new_n982_), .O(new_n1221_));
  AND      g1205(.a(new_n1221_), .b(new_n565_), .O(new_n1222_));
  AND      g1206(.a(new_n1222_), .b(new_n1220_), .O(new_n1223_));
  OR       g1207(.a(new_n1223_), .b(new_n1219_), .O(new_n1224_));
  AND      g1208(.a(new_n1224_), .b(new_n53_), .O(new_n1225_));
  OR       g1209(.a(i_2_3_99_0), .b(new_n53_), .O(new_n1226_));
  AND      g1210(.a(new_n742_), .b(new_n171_), .O(new_n1227_));
  AND      g1211(.a(new_n1227_), .b(new_n1226_), .O(new_n1228_));
  AND      g1212(.a(new_n206_), .b(new_n245_), .O(new_n1229_));
  OR       g1213(.a(new_n1229_), .b(new_n1228_), .O(new_n1230_));
  AND      g1214(.a(new_n1230_), .b(i_2_3_72_0), .O(new_n1231_));
  OR       g1215(.a(new_n952_), .b(new_n21_), .O(new_n1232_));
  AND      g1216(.a(new_n348_), .b(new_n278_), .O(new_n1233_));
  AND      g1217(.a(new_n1233_), .b(new_n1232_), .O(new_n1234_));
  OR       g1218(.a(new_n1234_), .b(new_n1231_), .O(new_n1235_));
  AND      g1219(.a(new_n1235_), .b(new_n18_), .O(new_n1236_));
  AND      g1220(.a(new_n462_), .b(new_n245_), .O(new_n1237_));
  OR       g1221(.a(new_n1237_), .b(new_n1236_), .O(new_n1238_));
  AND      g1222(.a(new_n1238_), .b(new_n688_), .O(new_n1239_));
  NOT      g1223(.a(new_n588_), .O(new_n1240_));
  AND      g1224(.a(new_n791_), .b(new_n1240_), .O(new_n1241_));
  OR       g1225(.a(new_n1241_), .b(new_n1239_), .O(new_n1242_));
  AND      g1226(.a(new_n1242_), .b(new_n105_), .O(new_n1243_));
  OR       g1227(.a(i_2_3_143_0), .b(new_n40_), .O(new_n1244_));
  AND      g1228(.a(new_n1244_), .b(new_n793_), .O(new_n1245_));
  OR       g1229(.a(new_n1245_), .b(i_2_3_43_0), .O(new_n1246_));
  NOT      g1230(.a(new_n893_), .O(new_n1247_));
  NAND     g1231(.a(new_n777_), .b(i_2_3_68_0), .O(new_n1248_));
  AND      g1232(.a(new_n1248_), .b(new_n1247_), .O(new_n1249_));
  AND      g1233(.a(new_n1249_), .b(new_n1246_), .O(new_n1250_));
  AND      g1234(.a(new_n1244_), .b(new_n480_), .O(new_n1251_));
  OR       g1235(.a(new_n1251_), .b(new_n1248_), .O(new_n1252_));
  AND      g1236(.a(new_n1252_), .b(i_2_3_79_0), .O(new_n1253_));
  OR       g1237(.a(new_n1253_), .b(i_2_3_77_0), .O(new_n1254_));
  OR       g1238(.a(new_n1254_), .b(new_n1250_), .O(new_n1255_));
  OR       g1239(.a(new_n908_), .b(i_2_3_68_0), .O(new_n1256_));
  AND      g1240(.a(new_n937_), .b(new_n780_), .O(new_n1257_));
  NAND     g1241(.a(new_n1257_), .b(new_n1256_), .O(new_n1258_));
  NAND     g1242(.a(new_n1258_), .b(new_n1255_), .O(new_n1259_));
  AND      g1243(.a(new_n1259_), .b(i_2_3_55_0), .O(new_n1260_));
  OR       g1244(.a(new_n846_), .b(new_n253_), .O(new_n1261_));
  NAND     g1245(.a(new_n1261_), .b(new_n512_), .O(new_n1262_));
  OR       g1246(.a(new_n1262_), .b(new_n697_), .O(new_n1263_));
  OR       g1247(.a(new_n1203_), .b(new_n30_), .O(new_n1264_));
  AND      g1248(.a(new_n1264_), .b(new_n206_), .O(new_n1265_));
  OR       g1249(.a(new_n1265_), .b(new_n756_), .O(new_n1266_));
  OR       g1250(.a(new_n1266_), .b(new_n1263_), .O(new_n1267_));
  AND      g1251(.a(new_n1267_), .b(new_n19_), .O(new_n1268_));
  NAND     g1252(.a(new_n1248_), .b(i_2_3_79_0), .O(new_n1269_));
  AND      g1253(.a(new_n1269_), .b(new_n756_), .O(new_n1270_));
  NAND     g1254(.a(new_n591_), .b(i_2_3_79_0), .O(new_n1271_));
  OR       g1255(.a(new_n1065_), .b(new_n212_), .O(new_n1272_));
  AND      g1256(.a(new_n1272_), .b(new_n928_), .O(new_n1273_));
  AND      g1257(.a(new_n1273_), .b(new_n1271_), .O(new_n1274_));
  OR       g1258(.a(new_n1274_), .b(new_n1270_), .O(new_n1275_));
  AND      g1259(.a(new_n1275_), .b(i_2_3_72_0), .O(new_n1276_));
  AND      g1260(.a(new_n597_), .b(new_n200_), .O(new_n1277_));
  AND      g1261(.a(new_n1277_), .b(new_n1256_), .O(new_n1278_));
  OR       g1262(.a(new_n1278_), .b(new_n1276_), .O(new_n1279_));
  OR       g1263(.a(new_n1279_), .b(new_n1268_), .O(new_n1280_));
  AND      g1264(.a(new_n1280_), .b(i_2_3_86_0), .O(new_n1281_));
  OR       g1265(.a(new_n1281_), .b(new_n1260_), .O(new_n1282_));
  AND      g1266(.a(new_n1282_), .b(new_n53_), .O(new_n1283_));
  OR       g1267(.a(new_n774_), .b(new_n721_), .O(new_n1284_));
  AND      g1268(.a(new_n1284_), .b(new_n77_), .O(new_n1285_));
  OR       g1269(.a(new_n1031_), .b(new_n886_), .O(new_n1286_));
  AND      g1270(.a(new_n1286_), .b(new_n21_), .O(new_n1287_));
  OR       g1271(.a(new_n1287_), .b(new_n1285_), .O(new_n1288_));
  AND      g1272(.a(new_n1288_), .b(new_n18_), .O(new_n1289_));
  AND      g1273(.a(new_n692_), .b(new_n511_), .O(new_n1290_));
  OR       g1274(.a(new_n1290_), .b(new_n1289_), .O(new_n1291_));
  AND      g1275(.a(new_n1291_), .b(new_n56_), .O(new_n1292_));
  NAND     g1276(.a(new_n252_), .b(new_n100_), .O(new_n1293_));
  AND      g1277(.a(new_n1293_), .b(new_n1154_), .O(new_n1294_));
  OR       g1278(.a(new_n1294_), .b(new_n1292_), .O(new_n1295_));
  OR       g1279(.a(new_n1295_), .b(new_n1283_), .O(new_n1296_));
  AND      g1280(.a(new_n1296_), .b(i_2_3_29_0), .O(new_n1297_));
  AND      g1281(.a(new_n688_), .b(new_n253_), .O(new_n1298_));
  AND      g1282(.a(new_n458_), .b(i_2_3_43_0), .O(new_n1299_));
  OR       g1283(.a(new_n1299_), .b(new_n1298_), .O(new_n1300_));
  AND      g1284(.a(new_n1300_), .b(i_2_3_72_0), .O(new_n1301_));
  AND      g1285(.a(new_n1000_), .b(new_n564_), .O(new_n1302_));
  OR       g1286(.a(new_n1302_), .b(new_n1301_), .O(new_n1303_));
  AND      g1287(.a(new_n1303_), .b(new_n53_), .O(new_n1304_));
  AND      g1288(.a(new_n772_), .b(new_n564_), .O(new_n1305_));
  OR       g1289(.a(new_n1305_), .b(new_n1304_), .O(new_n1306_));
  AND      g1290(.a(new_n1306_), .b(new_n18_), .O(new_n1307_));
  AND      g1291(.a(new_n739_), .b(new_n25_), .O(new_n1308_));
  AND      g1292(.a(new_n1308_), .b(new_n840_), .O(new_n1309_));
  OR       g1293(.a(new_n1309_), .b(new_n1307_), .O(new_n1310_));
  AND      g1294(.a(new_n1310_), .b(i_2_3_86_0), .O(new_n1311_));
  NOT      g1295(.a(new_n456_), .O(new_n1312_));
  AND      g1296(.a(new_n1154_), .b(new_n1312_), .O(new_n1313_));
  OR       g1297(.a(new_n1313_), .b(new_n1311_), .O(new_n1314_));
  AND      g1298(.a(new_n1314_), .b(new_n21_), .O(new_n1315_));
  AND      g1299(.a(new_n1019_), .b(new_n56_), .O(new_n1316_));
  AND      g1300(.a(new_n1316_), .b(new_n828_), .O(new_n1317_));
  OR       g1301(.a(new_n1317_), .b(new_n1315_), .O(new_n1318_));
  OR       g1302(.a(new_n1318_), .b(new_n1297_), .O(new_n1319_));
  AND      g1303(.a(new_n1319_), .b(new_n20_), .O(new_n1320_));
  OR       g1304(.a(new_n1320_), .b(new_n1243_), .O(new_n1321_));
  AND      g1305(.a(new_n1321_), .b(new_n31_), .O(new_n1322_));
  NOT      g1306(.a(new_n166_), .O(new_n1323_));
  AND      g1307(.a(new_n892_), .b(new_n1323_), .O(new_n1324_));
  AND      g1308(.a(new_n1324_), .b(new_n921_), .O(new_n1325_));
  OR       g1309(.a(new_n1325_), .b(new_n1322_), .O(new_n1326_));
  OR       g1310(.a(new_n1326_), .b(new_n1225_), .O(new_n1327_));
  OR       g1311(.a(new_n1327_), .b(new_n1192_), .O(new_n1328_));
  OR       g1312(.a(new_n1328_), .b(new_n873_), .O(o_2_3_0_0));
endmodule


